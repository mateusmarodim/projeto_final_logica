-- system_0.vhd

-- Generated using ACDS version 13.0sp1 232 at 2024.07.05.04:12:32

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_0 is
	port (
		clk_50                               : in    std_logic                     := '0';             --                   clk_50_clk_in.clk
		bidir_port_to_and_from_the_SD_DAT    : inout std_logic                     := '0';             --      SD_DAT_external_connection.export
		out_port_from_the_led_red            : out   std_logic_vector(17 downto 0);                    --     led_red_external_connection.export
		zs_addr_from_the_sdram_0             : out   std_logic_vector(11 downto 0);                    --                    sdram_0_wire.addr
		zs_ba_from_the_sdram_0               : out   std_logic_vector(1 downto 0);                     --                                .ba
		zs_cas_n_from_the_sdram_0            : out   std_logic;                                        --                                .cas_n
		zs_cke_from_the_sdram_0              : out   std_logic;                                        --                                .cke
		zs_cs_n_from_the_sdram_0             : out   std_logic;                                        --                                .cs_n
		zs_dq_to_and_from_the_sdram_0        : inout std_logic_vector(15 downto 0) := (others => '0'); --                                .dq
		zs_dqm_from_the_sdram_0              : out   std_logic_vector(1 downto 0);                     --                                .dqm
		zs_ras_n_from_the_sdram_0            : out   std_logic;                                        --                                .ras_n
		zs_we_n_from_the_sdram_0             : out   std_logic;                                        --                                .we_n
		tri_state_bridge_0_data              : inout std_logic_vector(7 downto 0)  := (others => '0'); -- tri_state_bridge_0_bridge_0_out.tri_state_bridge_0_data
		tri_state_bridge_0_readn             : out   std_logic_vector(0 downto 0);                     --                                .tri_state_bridge_0_readn
		write_n_to_the_cfi_flash_0           : out   std_logic_vector(0 downto 0);                     --                                .write_n_to_the_cfi_flash_0
		tri_state_bridge_0_address           : out   std_logic_vector(21 downto 0);                    --                                .tri_state_bridge_0_address
		select_n_to_the_cfi_flash_0          : out   std_logic_vector(0 downto 0);                     --                                .select_n_to_the_cfi_flash_0
		reset_n                              : in    std_logic                     := '0';             --          merged_resets_in_reset.reset_n
		bidir_port_to_and_from_the_SD_CMD    : inout std_logic                     := '0';             --      SD_CMD_external_connection.export
		in_port_to_the_button_pio            : in    std_logic_vector(3 downto 0)  := (others => '0'); --  button_pio_external_connection.export
		USB_DATA_to_and_from_the_ISP1362     : inout std_logic_vector(15 downto 0) := (others => '0'); --             ISP1362_conduit_end.DATA
		USB_ADDR_from_the_ISP1362            : out   std_logic_vector(1 downto 0);                     --                                .ADDR
		USB_RD_N_from_the_ISP1362            : out   std_logic;                                        --                                .RD_N
		USB_WR_N_from_the_ISP1362            : out   std_logic;                                        --                                .WR_N
		USB_CS_N_from_the_ISP1362            : out   std_logic;                                        --                                .CS_N
		USB_RST_N_from_the_ISP1362           : out   std_logic;                                        --                                .RST_N
		USB_INT0_to_the_ISP1362              : in    std_logic                     := '0';             --                                .INT0
		USB_INT1_to_the_ISP1362              : in    std_logic                     := '0';             --                                .INT1
		out_port_from_the_SD_CLK             : out   std_logic;                                        --      SD_CLK_external_connection.export
		out_port_from_the_led_green          : out   std_logic_vector(8 downto 0);                     --   led_green_external_connection.export
		in_port_to_the_switch_pio            : in    std_logic_vector(17 downto 0) := (others => '0'); --  switch_pio_external_connection.export
		LCD_RS_from_the_lcd_16207_0          : out   std_logic;                                        --            lcd_16207_0_external.RS
		LCD_RW_from_the_lcd_16207_0          : out   std_logic;                                        --                                .RW
		LCD_data_to_and_from_the_lcd_16207_0 : inout std_logic_vector(7 downto 0)  := (others => '0'); --                                .data
		LCD_E_from_the_lcd_16207_0           : out   std_logic;                                        --                                .E
		rxd_to_the_uart_0                    : in    std_logic                     := '0';             --      uart_0_external_connection.rxd
		txd_from_the_uart_0                  : out   std_logic;                                        --                                .txd
		audio_0_oAUD_DATA                    : out   std_logic;                                        --                         audio_0.oAUD_DATA
		audio_0_oAUD_LRCK                    : out   std_logic;                                        --                                .oAUD_LRCK
		audio_0_oAUD_BCK                     : out   std_logic;                                        --                                .oAUD_BCK
		audio_0_oAUD_XCK                     : out   std_logic;                                        --                                .oAUD_XCK
		audio_0_iCLK_18_4                    : in    std_logic                     := '0';             --                                .iCLK_18_4
		vga_0_VGA_R                          : out   std_logic_vector(9 downto 0);                     --                           vga_0.VGA_R
		vga_0_VGA_G                          : out   std_logic_vector(9 downto 0);                     --                                .VGA_G
		vga_0_VGA_B                          : out   std_logic_vector(9 downto 0);                     --                                .VGA_B
		vga_0_VGA_HS                         : out   std_logic;                                        --                                .VGA_HS
		vga_0_VGA_VS                         : out   std_logic;                                        --                                .VGA_VS
		vga_0_VGA_SYNC                       : out   std_logic;                                        --                                .VGA_SYNC
		vga_0_VGA_BLANK                      : out   std_logic;                                        --                                .VGA_BLANK
		vga_0_VGA_CLK                        : out   std_logic;                                        --                                .VGA_CLK
		vga_0_iCLK_25                        : in    std_logic                     := '0';             --                                .iCLK_25
		dm9000a_iOSC_50                      : in    std_logic                     := '0';             --                         dm9000a.iOSC_50
		dm9000a_ENET_DATA                    : inout std_logic_vector(15 downto 0) := (others => '0'); --                                .ENET_DATA
		dm9000a_ENET_CMD                     : out   std_logic;                                        --                                .ENET_CMD
		dm9000a_ENET_RD_N                    : out   std_logic;                                        --                                .ENET_RD_N
		dm9000a_ENET_WR_N                    : out   std_logic;                                        --                                .ENET_WR_N
		dm9000a_ENET_CS_N                    : out   std_logic;                                        --                                .ENET_CS_N
		dm9000a_ENET_RST_N                   : out   std_logic;                                        --                                .ENET_RST_N
		dm9000a_ENET_CLK                     : out   std_logic;                                        --                                .ENET_CLK
		dm9000a_ENET_INT                     : in    std_logic                     := '0';             --                                .ENET_INT
		seg7_display_oSEG0                   : out   std_logic_vector(6 downto 0);                     --                    seg7_display.oSEG0
		seg7_display_oSEG1                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG1
		seg7_display_oSEG2                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG2
		seg7_display_oSEG3                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG3
		seg7_display_oSEG4                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG4
		seg7_display_oSEG5                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG5
		seg7_display_oSEG6                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG6
		seg7_display_oSEG7                   : out   std_logic_vector(6 downto 0);                     --                                .oSEG7
		sram_0_avalon_slave_0_export_DQ      : inout std_logic_vector(15 downto 0) := (others => '0'); --    sram_0_avalon_slave_0_export.DQ
		sram_0_avalon_slave_0_export_ADDR    : out   std_logic_vector(17 downto 0);                    --                                .ADDR
		sram_0_avalon_slave_0_export_UB_N    : out   std_logic;                                        --                                .UB_N
		sram_0_avalon_slave_0_export_LB_N    : out   std_logic;                                        --                                .LB_N
		sram_0_avalon_slave_0_export_WE_N    : out   std_logic;                                        --                                .WE_N
		sram_0_avalon_slave_0_export_CE_N    : out   std_logic;                                        --                                .CE_N
		sram_0_avalon_slave_0_export_OE_N    : out   std_logic;                                        --                                .OE_N
		cw_output_export                     : out   std_logic;                                        --                       cw_output.export
		ccw_output_export                    : out   std_logic                                         --                      ccw_output.export
	);
end entity system_0;

architecture rtl of system_0 is
	component system_0_sdram_0 is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component system_0_sdram_0;

	component system_0_epcs_controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			dataavailable : out std_logic;                                        -- dataavailable
			endofpacket   : out std_logic;                                        -- endofpacket
			read_n        : in  std_logic                     := 'X';             -- read_n
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			readyfordata  : out std_logic;                                        -- readyfordata
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq           : out std_logic                                         -- irq
		);
	end component system_0_epcs_controller;

	component system_0_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component system_0_jtag_uart_0;

	component system_0_uart_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component system_0_uart_0;

	component system_0_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component system_0_timer_0;

	component system_0_lcd_16207_0 is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			LCD_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component system_0_lcd_16207_0;

	component system_0_led_red is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(17 downto 0)                     -- export
		);
	end component system_0_led_red;

	component system_0_led_green is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(8 downto 0)                      -- export
		);
	end component system_0_led_green;

	component system_0_button_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component system_0_button_pio;

	component system_0_switch_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(17 downto 0) := (others => 'X')  -- export
		);
	end component system_0_switch_pio;

	component system_0_SD_DAT is
		port (
			clk        : in    std_logic                     := 'X';             -- clk
			reset_n    : in    std_logic                     := 'X';             -- reset_n
			address    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in    std_logic                     := 'X';             -- write_n
			writedata  : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in    std_logic                     := 'X';             -- chipselect
			readdata   : out   std_logic_vector(31 downto 0);                    -- readdata
			bidir_port : inout std_logic                     := 'X'              -- export
		);
	end component system_0_SD_DAT;

	component system_0_SD_CLK is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component system_0_SD_CLK;

	component ISP1362_IF is
		port (
			avs_hc_clk_iCLK           : in    std_logic                     := 'X';             -- clk
			avs_hc_reset_n_iRST_N     : in    std_logic                     := 'X';             -- reset_n
			avs_hc_writedata_iDATA    : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_hc_readdata_oDATA     : out   std_logic_vector(15 downto 0);                    -- readdata
			avs_hc_address_iADDR      : in    std_logic                     := 'X';             -- address
			avs_hc_read_n_iRD_N       : in    std_logic                     := 'X';             -- read_n
			avs_hc_write_n_iWR_N      : in    std_logic                     := 'X';             -- write_n
			avs_hc_chipselect_n_iCS_N : in    std_logic                     := 'X';             -- chipselect_n
			avs_hc_irq_n_oINT0_N      : out   std_logic;                                        -- irq_n
			avs_dc_clk_iCLK           : in    std_logic                     := 'X';             -- clk
			avs_dc_reset_n_iRST_N     : in    std_logic                     := 'X';             -- reset_n
			avs_dc_writedata_iDATA    : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			avs_dc_readdata_oDATA     : out   std_logic_vector(15 downto 0);                    -- readdata
			avs_dc_address_iADDR      : in    std_logic                     := 'X';             -- address
			avs_dc_read_n_iRD_N       : in    std_logic                     := 'X';             -- read_n
			avs_dc_write_n_iWR_N      : in    std_logic                     := 'X';             -- write_n
			avs_dc_chipselect_n_iCS_N : in    std_logic                     := 'X';             -- chipselect_n
			avs_dc_irq_n_oINT0_N      : out   std_logic;                                        -- irq_n
			USB_DATA                  : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			USB_ADDR                  : out   std_logic_vector(1 downto 0);                     -- export
			USB_RD_N                  : out   std_logic;                                        -- export
			USB_WR_N                  : out   std_logic;                                        -- export
			USB_CS_N                  : out   std_logic;                                        -- export
			USB_RST_N                 : out   std_logic;                                        -- export
			USB_INT0                  : in    std_logic                     := 'X';             -- export
			USB_INT1                  : in    std_logic                     := 'X'              -- export
		);
	end component ISP1362_IF;

	component system_0_cpu_0 is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			d_address                             : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(24 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component system_0_cpu_0;

	component system_0_tri_state_bridge_0_bridge_0 is
		port (
			clk                               : in    std_logic                     := 'X';             -- clk
			reset                             : in    std_logic                     := 'X';             -- reset
			request                           : in    std_logic                     := 'X';             -- request
			grant                             : out   std_logic;                                        -- grant
			tcs_tri_state_bridge_0_data       : in    std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data_out
			tcs_tri_state_bridge_0_data_outen : in    std_logic                     := 'X';             -- tri_state_bridge_0_data_outen
			tcs_tri_state_bridge_0_data_in    : out   std_logic_vector(7 downto 0);                     -- tri_state_bridge_0_data_in
			tcs_tri_state_bridge_0_readn      : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- tri_state_bridge_0_readn_out
			tcs_write_n_to_the_cfi_flash_0    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_to_the_cfi_flash_0_out
			tcs_tri_state_bridge_0_address    : in    std_logic_vector(21 downto 0) := (others => 'X'); -- tri_state_bridge_0_address_out
			tcs_select_n_to_the_cfi_flash_0   : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- select_n_to_the_cfi_flash_0_out
			tri_state_bridge_0_data           : inout std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data
			tri_state_bridge_0_readn          : out   std_logic_vector(0 downto 0);                     -- tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0        : out   std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address        : out   std_logic_vector(21 downto 0);                    -- tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0       : out   std_logic_vector(0 downto 0)                      -- select_n_to_the_cfi_flash_0
		);
	end component system_0_tri_state_bridge_0_bridge_0;

	component system_0_tri_state_bridge_0_pinSharer_0 is
		port (
			clk_clk                       : in  std_logic                     := 'X';             -- clk
			reset_reset                   : in  std_logic                     := 'X';             -- reset
			request                       : out std_logic;                                        -- request
			grant                         : in  std_logic                     := 'X';             -- grant
			tri_state_bridge_0_address    : out std_logic_vector(21 downto 0);                    -- tri_state_bridge_0_address_out
			tri_state_bridge_0_readn      : out std_logic_vector(0 downto 0);                     -- tri_state_bridge_0_readn_out
			write_n_to_the_cfi_flash_0    : out std_logic_vector(0 downto 0);                     -- write_n_to_the_cfi_flash_0_out
			tri_state_bridge_0_data       : out std_logic_vector(7 downto 0);                     -- tri_state_bridge_0_data_out
			tri_state_bridge_0_data_in    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- tri_state_bridge_0_data_in
			tri_state_bridge_0_data_outen : out std_logic;                                        -- tri_state_bridge_0_data_outen
			select_n_to_the_cfi_flash_0   : out std_logic_vector(0 downto 0);                     -- select_n_to_the_cfi_flash_0_out
			tcs0_request                  : in  std_logic                     := 'X';             -- request
			tcs0_grant                    : out std_logic;                                        -- grant
			tcs0_address_out              : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address_out
			tcs0_read_n_out               : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- read_n_out
			tcs0_write_n_out              : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs0_data_out                 : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data_out
			tcs0_data_in                  : out std_logic_vector(7 downto 0);                     -- data_in
			tcs0_data_outen               : in  std_logic                     := 'X';             -- data_outen
			tcs0_chipselect_n_out         : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- chipselect_n_out
		);
	end component system_0_tri_state_bridge_0_pinSharer_0;

	component system_0_cfi_flash_0 is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			reset_reset          : in  std_logic                     := 'X';             -- reset
			uas_address          : in  std_logic_vector(21 downto 0) := (others => 'X'); -- address
			uas_burstcount       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uas_read             : in  std_logic                     := 'X';             -- read
			uas_write            : in  std_logic                     := 'X';             -- write
			uas_waitrequest      : out std_logic;                                        -- waitrequest
			uas_readdatavalid    : out std_logic;                                        -- readdatavalid
			uas_byteenable       : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata         : out std_logic_vector(7 downto 0);                     -- readdata
			uas_writedata        : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uas_lock             : in  std_logic                     := 'X';             -- lock
			uas_debugaccess      : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out      : out std_logic;                                        -- write_n_out
			tcm_read_n_out       : out std_logic;                                        -- read_n_out
			tcm_chipselect_n_out : out std_logic;                                        -- chipselect_n_out
			tcm_request          : out std_logic;                                        -- request
			tcm_grant            : in  std_logic                     := 'X';             -- grant
			tcm_address_out      : out std_logic_vector(21 downto 0);                    -- address_out
			tcm_data_out         : out std_logic_vector(7 downto 0);                     -- data_out
			tcm_data_outen       : out std_logic;                                        -- data_outen
			tcm_data_in          : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- data_in
		);
	end component system_0_cfi_flash_0;

	component system_0_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component system_0_sysid_qsys_0;

	component AUDIO_DAC_FIFO is
		generic (
			REF_CLK     : integer := 18432000;
			SAMPLE_RATE : integer := 48000;
			DATA_WIDTH  : integer := 16;
			CHANNEL_NUM : integer := 2
		);
		port (
			iWR_CLK   : in  std_logic                     := 'X';             -- clk
			iRST_N    : in  std_logic                     := 'X';             -- reset_n
			oAUD_DATA : out std_logic;                                        -- export
			oAUD_LRCK : out std_logic;                                        -- export
			oAUD_BCK  : out std_logic;                                        -- export
			oAUD_XCK  : out std_logic;                                        -- export
			iCLK_18_4 : in  std_logic                     := 'X';             -- export
			iDATA     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			iWR       : in  std_logic                     := 'X';             -- write
			oDATA     : out std_logic_vector(15 downto 0)                     -- readdata
		);
	end component AUDIO_DAC_FIFO;

	component VGA_NIOS_CTRL is
		generic (
			RAM_SIZE : integer := 307200
		);
		port (
			iCLK      : in  std_logic                     := 'X';             -- clk
			iRST_N    : in  std_logic                     := 'X';             -- reset_n
			VGA_R     : out std_logic_vector(9 downto 0);                     -- export
			VGA_G     : out std_logic_vector(9 downto 0);                     -- export
			VGA_B     : out std_logic_vector(9 downto 0);                     -- export
			VGA_HS    : out std_logic;                                        -- export
			VGA_VS    : out std_logic;                                        -- export
			VGA_SYNC  : out std_logic;                                        -- export
			VGA_BLANK : out std_logic;                                        -- export
			VGA_CLK   : out std_logic;                                        -- export
			iCLK_25   : in  std_logic                     := 'X';             -- export
			oDATA     : out std_logic_vector(15 downto 0);                    -- readdata
			iDATA     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			iADDR     : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			iWR       : in  std_logic                     := 'X';             -- write
			iRD       : in  std_logic                     := 'X';             -- read
			iCS       : in  std_logic                     := 'X'              -- chipselect
		);
	end component VGA_NIOS_CTRL;

	component DM9000A_IF is
		port (
			iCLK       : in    std_logic                     := 'X';             -- clk
			iRST_N     : in    std_logic                     := 'X';             -- reset_n
			iOSC_50    : in    std_logic                     := 'X';             -- export
			ENET_DATA  : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			ENET_CMD   : out   std_logic;                                        -- export
			ENET_RD_N  : out   std_logic;                                        -- export
			ENET_WR_N  : out   std_logic;                                        -- export
			ENET_CS_N  : out   std_logic;                                        -- export
			ENET_RST_N : out   std_logic;                                        -- export
			ENET_CLK   : out   std_logic;                                        -- export
			ENET_INT   : in    std_logic                     := 'X';             -- export
			iDATA      : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			iCMD       : in    std_logic                     := 'X';             -- address
			iRD_N      : in    std_logic                     := 'X';             -- read_n
			iWR_N      : in    std_logic                     := 'X';             -- write_n
			iCS_N      : in    std_logic                     := 'X';             -- chipselect_n
			oDATA      : out   std_logic_vector(15 downto 0);                    -- readdata
			oINT       : out   std_logic                                         -- irq
		);
	end component DM9000A_IF;

	component SEG7_LUT_8 is
		port (
			iCLK   : in  std_logic                     := 'X';             -- clk
			iRST_N : in  std_logic                     := 'X';             -- reset_n
			oSEG0  : out std_logic_vector(6 downto 0);                     -- export
			oSEG1  : out std_logic_vector(6 downto 0);                     -- export
			oSEG2  : out std_logic_vector(6 downto 0);                     -- export
			oSEG3  : out std_logic_vector(6 downto 0);                     -- export
			oSEG4  : out std_logic_vector(6 downto 0);                     -- export
			oSEG5  : out std_logic_vector(6 downto 0);                     -- export
			oSEG6  : out std_logic_vector(6 downto 0);                     -- export
			oSEG7  : out std_logic_vector(6 downto 0);                     -- export
			iDIG   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			iWR    : in  std_logic                     := 'X'              -- write
		);
	end component SEG7_LUT_8;

	component SRAM_16Bit_512K is
		port (
			iCLK      : in    std_logic                     := 'X';             -- clk
			iRST_N    : in    std_logic                     := 'X';             -- reset_n
			SRAM_DQ   : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			SRAM_ADDR : out   std_logic_vector(17 downto 0);                    -- export
			SRAM_UB_N : out   std_logic;                                        -- export
			SRAM_LB_N : out   std_logic;                                        -- export
			SRAM_WE_N : out   std_logic;                                        -- export
			SRAM_CE_N : out   std_logic;                                        -- export
			SRAM_OE_N : out   std_logic;                                        -- export
			iDATA     : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			oDATA     : out   std_logic_vector(15 downto 0);                    -- readdata
			iADDR     : in    std_logic_vector(17 downto 0) := (others => 'X'); -- address
			iWE_N     : in    std_logic                     := 'X';             -- write_n
			iOE_N     : in    std_logic                     := 'X';             -- read_n
			iCE_N     : in    std_logic                     := 'X';             -- chipselect_n
			iBE_N     : in    std_logic_vector(1 downto 0)  := (others => 'X')  -- byteenable_n
		);
	end component SRAM_16Bit_512K;

	component top_avalon is
		port (
			chipselect : in  std_logic                     := 'X';             -- chipselect
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			add        : in  std_logic                     := 'X';             -- address
			write_en   : in  std_logic                     := 'X';             -- write
			read_en    : in  std_logic                     := 'X';             -- read
			clock      : in  std_logic                     := 'X';             -- clk
			resetn     : in  std_logic                     := 'X'              -- reset_n
		);
	end component top_avalon;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			av_address              : in  std_logic_vector(24 downto 0)  := (others => 'X'); -- address
			av_write                : in  std_logic                      := 'X';             -- write
			av_read                 : in  std_logic                      := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                     -- readdata
			av_waitrequest          : out std_logic;                                         -- waitrequest
			av_readdatavalid        : out std_logic;                                         -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)   := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)   := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                      := 'X';             -- debugaccess
			av_lock                 : in  std_logic                      := 'X';             -- lock
			cp_valid                : out std_logic;                                         -- valid
			cp_data                 : out std_logic_vector(101 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_endofpacket          : out std_logic;                                         -- endofpacket
			cp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : in  std_logic                      := 'X';             -- valid
			rp_data                 : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                         -- ready
			av_response             : out std_logic_vector(1 downto 0);                      -- response
			av_writeresponserequest : in  std_logic                      := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                          -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component system_0_addr_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component system_0_addr_router;

	component system_0_addr_router_001 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component system_0_addr_router_001;

	component system_0_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component system_0_id_router;

	component system_0_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(83 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component system_0_id_router_001;

	component system_0_id_router_003 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(74 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(74 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component system_0_id_router_003;

	component system_0_id_router_005 is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(101 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component system_0_id_router_005;

	component system_0_id_router_023 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(83 downto 0);                    -- data
			src_channel        : out std_logic_vector(26 downto 0);                    -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component system_0_id_router_023;

	component altera_merlin_traffic_limiter is
		generic (
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_TRANS_POSTED          : integer := 0;
			PKT_TRANS_WRITE           : integer := 0;
			MAX_OUTSTANDING_RESPONSES : integer := 0;
			PIPELINED                 : integer := 0;
			ST_DATA_W                 : integer := 72;
			ST_CHANNEL_W              : integer := 1;
			VALID_WIDTH               : integer := 1;
			ENFORCE_ORDER             : integer := 1;
			PREVENT_HAZARDS           : integer := 0;
			PKT_BYTE_CNT_H            : integer := 0;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 0;
			PKT_BYTEEN_L              : integer := 0
		);
		port (
			clk                    : in  std_logic                      := 'X';             -- clk
			reset                  : in  std_logic                      := 'X';             -- reset
			cmd_sink_ready         : out std_logic;                                         -- ready
			cmd_sink_valid         : in  std_logic                      := 'X';             -- valid
			cmd_sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			cmd_sink_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			cmd_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			cmd_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			cmd_src_ready          : in  std_logic                      := 'X';             -- ready
			cmd_src_data           : out std_logic_vector(101 downto 0);                    -- data
			cmd_src_channel        : out std_logic_vector(26 downto 0);                     -- channel
			cmd_src_startofpacket  : out std_logic;                                         -- startofpacket
			cmd_src_endofpacket    : out std_logic;                                         -- endofpacket
			rsp_sink_ready         : out std_logic;                                         -- ready
			rsp_sink_valid         : in  std_logic                      := 'X';             -- valid
			rsp_sink_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			rsp_sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			rsp_sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			rsp_sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			rsp_src_ready          : in  std_logic                      := 'X';             -- ready
			rsp_src_valid          : out std_logic;                                         -- valid
			rsp_src_data           : out std_logic_vector(101 downto 0);                    -- data
			rsp_src_channel        : out std_logic_vector(26 downto 0);                     -- channel
			rsp_src_startofpacket  : out std_logic;                                         -- startofpacket
			rsp_src_endofpacket    : out std_logic;                                         -- endofpacket
			cmd_src_valid          : out std_logic_vector(26 downto 0)                      -- data
		);
	end component altera_merlin_traffic_limiter;

	component system_0_cmd_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- data
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(101 downto 0);                    -- data
			src1_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic;                                         -- endofpacket
			src2_ready         : in  std_logic                      := 'X';             -- ready
			src2_valid         : out std_logic;                                         -- valid
			src2_data          : out std_logic_vector(101 downto 0);                    -- data
			src2_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src2_startofpacket : out std_logic;                                         -- startofpacket
			src2_endofpacket   : out std_logic;                                         -- endofpacket
			src3_ready         : in  std_logic                      := 'X';             -- ready
			src3_valid         : out std_logic;                                         -- valid
			src3_data          : out std_logic_vector(101 downto 0);                    -- data
			src3_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src3_startofpacket : out std_logic;                                         -- startofpacket
			src3_endofpacket   : out std_logic;                                         -- endofpacket
			src4_ready         : in  std_logic                      := 'X';             -- ready
			src4_valid         : out std_logic;                                         -- valid
			src4_data          : out std_logic_vector(101 downto 0);                    -- data
			src4_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src4_startofpacket : out std_logic;                                         -- startofpacket
			src4_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component system_0_cmd_xbar_demux;

	component system_0_cmd_xbar_demux_001 is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			sink_ready          : out std_logic;                                         -- ready
			sink_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink_valid          : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready          : in  std_logic                      := 'X';             -- ready
			src0_valid          : out std_logic;                                         -- valid
			src0_data           : out std_logic_vector(101 downto 0);                    -- data
			src0_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src0_startofpacket  : out std_logic;                                         -- startofpacket
			src0_endofpacket    : out std_logic;                                         -- endofpacket
			src1_ready          : in  std_logic                      := 'X';             -- ready
			src1_valid          : out std_logic;                                         -- valid
			src1_data           : out std_logic_vector(101 downto 0);                    -- data
			src1_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src1_startofpacket  : out std_logic;                                         -- startofpacket
			src1_endofpacket    : out std_logic;                                         -- endofpacket
			src2_ready          : in  std_logic                      := 'X';             -- ready
			src2_valid          : out std_logic;                                         -- valid
			src2_data           : out std_logic_vector(101 downto 0);                    -- data
			src2_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src2_startofpacket  : out std_logic;                                         -- startofpacket
			src2_endofpacket    : out std_logic;                                         -- endofpacket
			src3_ready          : in  std_logic                      := 'X';             -- ready
			src3_valid          : out std_logic;                                         -- valid
			src3_data           : out std_logic_vector(101 downto 0);                    -- data
			src3_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src3_startofpacket  : out std_logic;                                         -- startofpacket
			src3_endofpacket    : out std_logic;                                         -- endofpacket
			src4_ready          : in  std_logic                      := 'X';             -- ready
			src4_valid          : out std_logic;                                         -- valid
			src4_data           : out std_logic_vector(101 downto 0);                    -- data
			src4_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src4_startofpacket  : out std_logic;                                         -- startofpacket
			src4_endofpacket    : out std_logic;                                         -- endofpacket
			src5_ready          : in  std_logic                      := 'X';             -- ready
			src5_valid          : out std_logic;                                         -- valid
			src5_data           : out std_logic_vector(101 downto 0);                    -- data
			src5_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src5_startofpacket  : out std_logic;                                         -- startofpacket
			src5_endofpacket    : out std_logic;                                         -- endofpacket
			src6_ready          : in  std_logic                      := 'X';             -- ready
			src6_valid          : out std_logic;                                         -- valid
			src6_data           : out std_logic_vector(101 downto 0);                    -- data
			src6_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src6_startofpacket  : out std_logic;                                         -- startofpacket
			src6_endofpacket    : out std_logic;                                         -- endofpacket
			src7_ready          : in  std_logic                      := 'X';             -- ready
			src7_valid          : out std_logic;                                         -- valid
			src7_data           : out std_logic_vector(101 downto 0);                    -- data
			src7_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src7_startofpacket  : out std_logic;                                         -- startofpacket
			src7_endofpacket    : out std_logic;                                         -- endofpacket
			src8_ready          : in  std_logic                      := 'X';             -- ready
			src8_valid          : out std_logic;                                         -- valid
			src8_data           : out std_logic_vector(101 downto 0);                    -- data
			src8_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src8_startofpacket  : out std_logic;                                         -- startofpacket
			src8_endofpacket    : out std_logic;                                         -- endofpacket
			src9_ready          : in  std_logic                      := 'X';             -- ready
			src9_valid          : out std_logic;                                         -- valid
			src9_data           : out std_logic_vector(101 downto 0);                    -- data
			src9_channel        : out std_logic_vector(26 downto 0);                     -- channel
			src9_startofpacket  : out std_logic;                                         -- startofpacket
			src9_endofpacket    : out std_logic;                                         -- endofpacket
			src10_ready         : in  std_logic                      := 'X';             -- ready
			src10_valid         : out std_logic;                                         -- valid
			src10_data          : out std_logic_vector(101 downto 0);                    -- data
			src10_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src10_startofpacket : out std_logic;                                         -- startofpacket
			src10_endofpacket   : out std_logic;                                         -- endofpacket
			src11_ready         : in  std_logic                      := 'X';             -- ready
			src11_valid         : out std_logic;                                         -- valid
			src11_data          : out std_logic_vector(101 downto 0);                    -- data
			src11_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src11_startofpacket : out std_logic;                                         -- startofpacket
			src11_endofpacket   : out std_logic;                                         -- endofpacket
			src12_ready         : in  std_logic                      := 'X';             -- ready
			src12_valid         : out std_logic;                                         -- valid
			src12_data          : out std_logic_vector(101 downto 0);                    -- data
			src12_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src12_startofpacket : out std_logic;                                         -- startofpacket
			src12_endofpacket   : out std_logic;                                         -- endofpacket
			src13_ready         : in  std_logic                      := 'X';             -- ready
			src13_valid         : out std_logic;                                         -- valid
			src13_data          : out std_logic_vector(101 downto 0);                    -- data
			src13_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src13_startofpacket : out std_logic;                                         -- startofpacket
			src13_endofpacket   : out std_logic;                                         -- endofpacket
			src14_ready         : in  std_logic                      := 'X';             -- ready
			src14_valid         : out std_logic;                                         -- valid
			src14_data          : out std_logic_vector(101 downto 0);                    -- data
			src14_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src14_startofpacket : out std_logic;                                         -- startofpacket
			src14_endofpacket   : out std_logic;                                         -- endofpacket
			src15_ready         : in  std_logic                      := 'X';             -- ready
			src15_valid         : out std_logic;                                         -- valid
			src15_data          : out std_logic_vector(101 downto 0);                    -- data
			src15_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src15_startofpacket : out std_logic;                                         -- startofpacket
			src15_endofpacket   : out std_logic;                                         -- endofpacket
			src16_ready         : in  std_logic                      := 'X';             -- ready
			src16_valid         : out std_logic;                                         -- valid
			src16_data          : out std_logic_vector(101 downto 0);                    -- data
			src16_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src16_startofpacket : out std_logic;                                         -- startofpacket
			src16_endofpacket   : out std_logic;                                         -- endofpacket
			src17_ready         : in  std_logic                      := 'X';             -- ready
			src17_valid         : out std_logic;                                         -- valid
			src17_data          : out std_logic_vector(101 downto 0);                    -- data
			src17_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src17_startofpacket : out std_logic;                                         -- startofpacket
			src17_endofpacket   : out std_logic;                                         -- endofpacket
			src18_ready         : in  std_logic                      := 'X';             -- ready
			src18_valid         : out std_logic;                                         -- valid
			src18_data          : out std_logic_vector(101 downto 0);                    -- data
			src18_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src18_startofpacket : out std_logic;                                         -- startofpacket
			src18_endofpacket   : out std_logic;                                         -- endofpacket
			src19_ready         : in  std_logic                      := 'X';             -- ready
			src19_valid         : out std_logic;                                         -- valid
			src19_data          : out std_logic_vector(101 downto 0);                    -- data
			src19_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src19_startofpacket : out std_logic;                                         -- startofpacket
			src19_endofpacket   : out std_logic;                                         -- endofpacket
			src20_ready         : in  std_logic                      := 'X';             -- ready
			src20_valid         : out std_logic;                                         -- valid
			src20_data          : out std_logic_vector(101 downto 0);                    -- data
			src20_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src20_startofpacket : out std_logic;                                         -- startofpacket
			src20_endofpacket   : out std_logic;                                         -- endofpacket
			src21_ready         : in  std_logic                      := 'X';             -- ready
			src21_valid         : out std_logic;                                         -- valid
			src21_data          : out std_logic_vector(101 downto 0);                    -- data
			src21_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src21_startofpacket : out std_logic;                                         -- startofpacket
			src21_endofpacket   : out std_logic;                                         -- endofpacket
			src22_ready         : in  std_logic                      := 'X';             -- ready
			src22_valid         : out std_logic;                                         -- valid
			src22_data          : out std_logic_vector(101 downto 0);                    -- data
			src22_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src22_startofpacket : out std_logic;                                         -- startofpacket
			src22_endofpacket   : out std_logic;                                         -- endofpacket
			src23_ready         : in  std_logic                      := 'X';             -- ready
			src23_valid         : out std_logic;                                         -- valid
			src23_data          : out std_logic_vector(101 downto 0);                    -- data
			src23_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src23_startofpacket : out std_logic;                                         -- startofpacket
			src23_endofpacket   : out std_logic;                                         -- endofpacket
			src24_ready         : in  std_logic                      := 'X';             -- ready
			src24_valid         : out std_logic;                                         -- valid
			src24_data          : out std_logic_vector(101 downto 0);                    -- data
			src24_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src24_startofpacket : out std_logic;                                         -- startofpacket
			src24_endofpacket   : out std_logic;                                         -- endofpacket
			src25_ready         : in  std_logic                      := 'X';             -- ready
			src25_valid         : out std_logic;                                         -- valid
			src25_data          : out std_logic_vector(101 downto 0);                    -- data
			src25_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src25_startofpacket : out std_logic;                                         -- startofpacket
			src25_endofpacket   : out std_logic;                                         -- endofpacket
			src26_ready         : in  std_logic                      := 'X';             -- ready
			src26_valid         : out std_logic;                                         -- valid
			src26_data          : out std_logic_vector(101 downto 0);                    -- data
			src26_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src26_startofpacket : out std_logic;                                         -- startofpacket
			src26_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component system_0_cmd_xbar_demux_001;

	component system_0_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(101 downto 0);                    -- data
			src_channel         : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component system_0_cmd_xbar_mux;

	component system_0_rsp_xbar_demux is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic;                                         -- endofpacket
			src1_ready         : in  std_logic                      := 'X';             -- ready
			src1_valid         : out std_logic;                                         -- valid
			src1_data          : out std_logic_vector(101 downto 0);                    -- data
			src1_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                         -- startofpacket
			src1_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component system_0_rsp_xbar_demux;

	component system_0_rsp_xbar_demux_005 is
		port (
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			sink_ready         : out std_logic;                                         -- ready
			sink_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)   := (others => 'X'); -- valid
			src0_ready         : in  std_logic                      := 'X';             -- ready
			src0_valid         : out std_logic;                                         -- valid
			src0_data          : out std_logic_vector(101 downto 0);                    -- data
			src0_channel       : out std_logic_vector(26 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                         -- startofpacket
			src0_endofpacket   : out std_logic                                          -- endofpacket
		);
	end component system_0_rsp_xbar_demux_005;

	component system_0_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                      := 'X';             -- clk
			reset               : in  std_logic                      := 'X';             -- reset
			src_ready           : in  std_logic                      := 'X';             -- ready
			src_valid           : out std_logic;                                         -- valid
			src_data            : out std_logic_vector(101 downto 0);                    -- data
			src_channel         : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                         -- startofpacket
			src_endofpacket     : out std_logic;                                         -- endofpacket
			sink0_ready         : out std_logic;                                         -- ready
			sink0_valid         : in  std_logic                      := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                         -- ready
			sink1_valid         : in  std_logic                      := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready         : out std_logic;                                         -- ready
			sink2_valid         : in  std_logic                      := 'X';             -- valid
			sink2_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink2_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink2_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready         : out std_logic;                                         -- ready
			sink3_valid         : in  std_logic                      := 'X';             -- valid
			sink3_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink3_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink3_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready         : out std_logic;                                         -- ready
			sink4_valid         : in  std_logic                      := 'X';             -- valid
			sink4_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink4_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink4_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component system_0_rsp_xbar_mux;

	component system_0_rsp_xbar_mux_001 is
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			src_ready            : in  std_logic                      := 'X';             -- ready
			src_valid            : out std_logic;                                         -- valid
			src_data             : out std_logic_vector(101 downto 0);                    -- data
			src_channel          : out std_logic_vector(26 downto 0);                     -- channel
			src_startofpacket    : out std_logic;                                         -- startofpacket
			src_endofpacket      : out std_logic;                                         -- endofpacket
			sink0_ready          : out std_logic;                                         -- ready
			sink0_valid          : in  std_logic                      := 'X';             -- valid
			sink0_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink0_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink0_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink0_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink1_ready          : out std_logic;                                         -- ready
			sink1_valid          : in  std_logic                      := 'X';             -- valid
			sink1_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink1_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink1_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink1_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink2_ready          : out std_logic;                                         -- ready
			sink2_valid          : in  std_logic                      := 'X';             -- valid
			sink2_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink2_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink2_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink2_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink3_ready          : out std_logic;                                         -- ready
			sink3_valid          : in  std_logic                      := 'X';             -- valid
			sink3_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink3_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink3_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink3_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink4_ready          : out std_logic;                                         -- ready
			sink4_valid          : in  std_logic                      := 'X';             -- valid
			sink4_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink4_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink4_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink4_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink5_ready          : out std_logic;                                         -- ready
			sink5_valid          : in  std_logic                      := 'X';             -- valid
			sink5_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink5_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink5_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink5_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink6_ready          : out std_logic;                                         -- ready
			sink6_valid          : in  std_logic                      := 'X';             -- valid
			sink6_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink6_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink6_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink6_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink7_ready          : out std_logic;                                         -- ready
			sink7_valid          : in  std_logic                      := 'X';             -- valid
			sink7_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink7_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink7_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink7_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink8_ready          : out std_logic;                                         -- ready
			sink8_valid          : in  std_logic                      := 'X';             -- valid
			sink8_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink8_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink8_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink8_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink9_ready          : out std_logic;                                         -- ready
			sink9_valid          : in  std_logic                      := 'X';             -- valid
			sink9_channel        : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink9_data           : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink9_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			sink9_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			sink10_ready         : out std_logic;                                         -- ready
			sink10_valid         : in  std_logic                      := 'X';             -- valid
			sink10_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink10_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink10_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink10_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink11_ready         : out std_logic;                                         -- ready
			sink11_valid         : in  std_logic                      := 'X';             -- valid
			sink11_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink11_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink11_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink11_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink12_ready         : out std_logic;                                         -- ready
			sink12_valid         : in  std_logic                      := 'X';             -- valid
			sink12_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink12_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink12_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink12_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink13_ready         : out std_logic;                                         -- ready
			sink13_valid         : in  std_logic                      := 'X';             -- valid
			sink13_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink13_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink13_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink13_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink14_ready         : out std_logic;                                         -- ready
			sink14_valid         : in  std_logic                      := 'X';             -- valid
			sink14_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink14_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink14_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink14_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink15_ready         : out std_logic;                                         -- ready
			sink15_valid         : in  std_logic                      := 'X';             -- valid
			sink15_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink15_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink15_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink15_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink16_ready         : out std_logic;                                         -- ready
			sink16_valid         : in  std_logic                      := 'X';             -- valid
			sink16_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink16_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink16_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink16_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink17_ready         : out std_logic;                                         -- ready
			sink17_valid         : in  std_logic                      := 'X';             -- valid
			sink17_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink17_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink17_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink17_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink18_ready         : out std_logic;                                         -- ready
			sink18_valid         : in  std_logic                      := 'X';             -- valid
			sink18_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink18_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink18_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink18_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink19_ready         : out std_logic;                                         -- ready
			sink19_valid         : in  std_logic                      := 'X';             -- valid
			sink19_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink19_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink19_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink19_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink20_ready         : out std_logic;                                         -- ready
			sink20_valid         : in  std_logic                      := 'X';             -- valid
			sink20_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink20_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink20_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink20_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink21_ready         : out std_logic;                                         -- ready
			sink21_valid         : in  std_logic                      := 'X';             -- valid
			sink21_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink21_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink21_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink21_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink22_ready         : out std_logic;                                         -- ready
			sink22_valid         : in  std_logic                      := 'X';             -- valid
			sink22_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink22_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink22_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink22_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink23_ready         : out std_logic;                                         -- ready
			sink23_valid         : in  std_logic                      := 'X';             -- valid
			sink23_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink23_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink23_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink23_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink24_ready         : out std_logic;                                         -- ready
			sink24_valid         : in  std_logic                      := 'X';             -- valid
			sink24_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink24_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink24_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink24_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink25_ready         : out std_logic;                                         -- ready
			sink25_valid         : in  std_logic                      := 'X';             -- valid
			sink25_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink25_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink25_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink25_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			sink26_ready         : out std_logic;                                         -- ready
			sink26_valid         : in  std_logic                      := 'X';             -- valid
			sink26_channel       : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			sink26_data          : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			sink26_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink26_endofpacket   : in  std_logic                      := 'X'              -- endofpacket
		);
	end component system_0_rsp_xbar_mux_001;

	component system_0_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			receiver4_irq : in  std_logic                     := 'X'; -- irq
			receiver5_irq : in  std_logic                     := 'X'; -- irq
			receiver6_irq : in  std_logic                     := 'X'; -- irq
			receiver7_irq : in  std_logic                     := 'X'; -- irq
			receiver8_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component system_0_irq_mapper;

	component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(102 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(102 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(84 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(84 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(17 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(75 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			out_data          : out std_logic_vector(9 downto 0);                     -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo;

	component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(101 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(102 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(102 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent;

	component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(1 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(1 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(15 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(83 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(26 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(84 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(84 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(17 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent;

	component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(24 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(0 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(0 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(7 downto 0);                     -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(74 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(74 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(26 downto 0) := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(75 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(75 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(9 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent;

	component system_0_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(83 downto 0);                     -- data
			out_channel          : out std_logic_vector(26 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component system_0_width_adapter;

	component system_0_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(83 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(101 downto 0);                    -- data
			out_channel          : out std_logic_vector(26 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component system_0_width_adapter_001;

	component system_0_width_adapter_002 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(101 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(74 downto 0);                     -- data
			out_channel          : out std_logic_vector(26 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component system_0_width_adapter_002;

	component system_0_width_adapter_003 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(26 downto 0)  := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(74 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(101 downto 0);                    -- data
			out_channel          : out std_logic_vector(26 downto 0);                     -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component system_0_width_adapter_003;

	component system_0_cpu_0_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component system_0_cpu_0_instruction_master_translator;

	component system_0_cpu_0_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(24 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component system_0_cpu_0_data_master_translator;

	component system_0_burst_adapter is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(26 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(83 downto 0);                    -- data
			source0_channel       : out std_logic_vector(26 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component system_0_burst_adapter;

	component system_0_burst_adapter_001 is
		generic (
			PKT_ADDR_H                : integer := 79;
			PKT_ADDR_L                : integer := 48;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BYTE_CNT_H            : integer := 5;
			PKT_BYTE_CNT_L            : integer := 0;
			PKT_BYTEEN_H              : integer := 83;
			PKT_BYTEEN_L              : integer := 80;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 88;
			PKT_BURST_TYPE_L          : integer := 87;
			PKT_BURSTWRAP_H           : integer := 11;
			PKT_BURSTWRAP_L           : integer := 6;
			PKT_TRANS_COMPRESSED_READ : integer := 14;
			PKT_TRANS_WRITE           : integer := 13;
			PKT_TRANS_READ            : integer := 12;
			OUT_NARROW_SIZE           : integer := 0;
			IN_NARROW_SIZE            : integer := 0;
			OUT_FIXED                 : integer := 0;
			OUT_COMPLETE_WRAP         : integer := 0;
			ST_DATA_W                 : integer := 89;
			ST_CHANNEL_W              : integer := 8;
			OUT_BYTE_CNT_H            : integer := 5;
			OUT_BURSTWRAP_H           : integer := 11;
			COMPRESSED_READ_SUPPORT   : integer := 1;
			BYTEENABLE_SYNTHESIS      : integer := 0;
			PIPE_INPUTS               : integer := 0;
			NO_WRAP_SUPPORT           : integer := 0;
			BURSTWRAP_CONST_MASK      : integer := 0;
			BURSTWRAP_CONST_VALUE     : integer := -1
		);
		port (
			clk                   : in  std_logic                     := 'X';             -- clk
			reset                 : in  std_logic                     := 'X';             -- reset
			sink0_valid           : in  std_logic                     := 'X';             -- valid
			sink0_data            : in  std_logic_vector(74 downto 0) := (others => 'X'); -- data
			sink0_channel         : in  std_logic_vector(26 downto 0) := (others => 'X'); -- channel
			sink0_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			sink0_ready           : out std_logic;                                        -- ready
			source0_valid         : out std_logic;                                        -- valid
			source0_data          : out std_logic_vector(74 downto 0);                    -- data
			source0_channel       : out std_logic_vector(26 downto 0);                    -- channel
			source0_startofpacket : out std_logic;                                        -- startofpacket
			source0_endofpacket   : out std_logic;                                        -- endofpacket
			source0_ready         : in  std_logic                     := 'X'              -- ready
		);
	end component system_0_burst_adapter_001;

	component system_0_cpu_0_jtag_debug_module_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_cpu_0_jtag_debug_module_translator;

	component system_0_sdram_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_sdram_0_s1_translator;

	component system_0_epcs_controller_epcs_control_port_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(8 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_epcs_controller_epcs_control_port_translator;

	component system_0_cfi_flash_0_uas_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(7 downto 0);                     -- readdata
			uav_writedata            : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(21 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_lock                  : out std_logic;                                        -- lock
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_cfi_flash_0_uas_translator;

	component system_0_sysid_qsys_0_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_sysid_qsys_0_control_slave_translator;

	component system_0_jtag_uart_0_avalon_jtag_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_jtag_uart_0_avalon_jtag_slave_translator;

	component system_0_uart_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_chipselect            : out std_logic;                                        -- chipselect
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_uart_0_s1_translator;

	component system_0_timer_0_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(2 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_timer_0_s1_translator;

	component system_0_lcd_16207_0_control_slave_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_lcd_16207_0_control_slave_translator;

	component system_0_led_red_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_led_red_s1_translator;

	component system_0_switch_pio_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(1 downto 0);                     -- address
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_switch_pio_s1_translator;

	component system_0_isp1362_hc_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_isp1362_hc_translator;

	component system_0_audio_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_audio_0_avalon_slave_0_translator;

	component system_0_vga_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(18 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_vga_0_avalon_slave_0_translator;

	component system_0_seg7_display_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_write                 : out std_logic;                                        -- write
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(0 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(0 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_seg7_display_avalon_slave_0_translator;

	component system_0_sram_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(15 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(17 downto 0);                    -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(15 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(1 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(1 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_sram_0_avalon_slave_0_translator;

	component system_0_lab7_final_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component system_0_lab7_final_0_avalon_slave_0_translator;

	component system_0_rst_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			reset_in1  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component system_0_rst_controller;

	component system_0_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component system_0_rst_controller_002;

	signal tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out                                     : std_logic_vector(0 downto 0);   -- tri_state_bridge_0_pinSharer_0:select_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_select_n_to_the_cfi_flash_0
	signal tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out                                      : std_logic_vector(21 downto 0);  -- tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_address -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_address
	signal tri_state_bridge_0_pinsharer_0_tcm_grant                                                               : std_logic;                      -- tri_state_bridge_0_bridge_0:grant -> tri_state_bridge_0_pinSharer_0:grant
	signal tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out                                        : std_logic_vector(0 downto 0);   -- tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_readn -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_readn
	signal tri_state_bridge_0_pinsharer_0_tcm_request                                                             : std_logic;                      -- tri_state_bridge_0_pinSharer_0:request -> tri_state_bridge_0_bridge_0:request
	signal tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in                                          : std_logic_vector(7 downto 0);   -- tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_in -> tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_in
	signal tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen                                       : std_logic;                      -- tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data_outen -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data_outen
	signal tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out                                      : std_logic_vector(0 downto 0);   -- tri_state_bridge_0_pinSharer_0:write_n_to_the_cfi_flash_0 -> tri_state_bridge_0_bridge_0:tcs_write_n_to_the_cfi_flash_0
	signal tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out                                         : std_logic_vector(7 downto 0);   -- tri_state_bridge_0_pinSharer_0:tri_state_bridge_0_data -> tri_state_bridge_0_bridge_0:tcs_tri_state_bridge_0_data
	signal cfi_flash_0_tcm_chipselect_n_out                                                                       : std_logic;                      -- cfi_flash_0:tcm_chipselect_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_chipselect_n_out
	signal cfi_flash_0_tcm_grant                                                                                  : std_logic;                      -- tri_state_bridge_0_pinSharer_0:tcs0_grant -> cfi_flash_0:tcm_grant
	signal cfi_flash_0_tcm_data_outen                                                                             : std_logic;                      -- cfi_flash_0:tcm_data_outen -> tri_state_bridge_0_pinSharer_0:tcs0_data_outen
	signal cfi_flash_0_tcm_request                                                                                : std_logic;                      -- cfi_flash_0:tcm_request -> tri_state_bridge_0_pinSharer_0:tcs0_request
	signal cfi_flash_0_tcm_data_out                                                                               : std_logic_vector(7 downto 0);   -- cfi_flash_0:tcm_data_out -> tri_state_bridge_0_pinSharer_0:tcs0_data_out
	signal cfi_flash_0_tcm_write_n_out                                                                            : std_logic;                      -- cfi_flash_0:tcm_write_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_write_n_out
	signal cfi_flash_0_tcm_address_out                                                                            : std_logic_vector(21 downto 0);  -- cfi_flash_0:tcm_address_out -> tri_state_bridge_0_pinSharer_0:tcs0_address_out
	signal cfi_flash_0_tcm_data_in                                                                                : std_logic_vector(7 downto 0);   -- tri_state_bridge_0_pinSharer_0:tcs0_data_in -> cfi_flash_0:tcm_data_in
	signal cfi_flash_0_tcm_read_n_out                                                                             : std_logic;                      -- cfi_flash_0:tcm_read_n_out -> tri_state_bridge_0_pinSharer_0:tcs0_read_n_out
	signal cpu_0_instruction_master_waitrequest                                                                   : std_logic;                      -- cpu_0_instruction_master_translator:av_waitrequest -> cpu_0:i_waitrequest
	signal cpu_0_instruction_master_address                                                                       : std_logic_vector(24 downto 0);  -- cpu_0:i_address -> cpu_0_instruction_master_translator:av_address
	signal cpu_0_instruction_master_read                                                                          : std_logic;                      -- cpu_0:i_read -> cpu_0_instruction_master_translator:av_read
	signal cpu_0_instruction_master_readdata                                                                      : std_logic_vector(31 downto 0);  -- cpu_0_instruction_master_translator:av_readdata -> cpu_0:i_readdata
	signal cpu_0_instruction_master_readdatavalid                                                                 : std_logic;                      -- cpu_0_instruction_master_translator:av_readdatavalid -> cpu_0:i_readdatavalid
	signal cpu_0_data_master_waitrequest                                                                          : std_logic;                      -- cpu_0_data_master_translator:av_waitrequest -> cpu_0:d_waitrequest
	signal cpu_0_data_master_writedata                                                                            : std_logic_vector(31 downto 0);  -- cpu_0:d_writedata -> cpu_0_data_master_translator:av_writedata
	signal cpu_0_data_master_address                                                                              : std_logic_vector(24 downto 0);  -- cpu_0:d_address -> cpu_0_data_master_translator:av_address
	signal cpu_0_data_master_write                                                                                : std_logic;                      -- cpu_0:d_write -> cpu_0_data_master_translator:av_write
	signal cpu_0_data_master_read                                                                                 : std_logic;                      -- cpu_0:d_read -> cpu_0_data_master_translator:av_read
	signal cpu_0_data_master_readdata                                                                             : std_logic_vector(31 downto 0);  -- cpu_0_data_master_translator:av_readdata -> cpu_0:d_readdata
	signal cpu_0_data_master_debugaccess                                                                          : std_logic;                      -- cpu_0:jtag_debug_module_debugaccess_to_roms -> cpu_0_data_master_translator:av_debugaccess
	signal cpu_0_data_master_byteenable                                                                           : std_logic_vector(3 downto 0);   -- cpu_0:d_byteenable -> cpu_0_data_master_translator:av_byteenable
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest                                     : std_logic;                      -- cpu_0:jtag_debug_module_waitrequest -> cpu_0_jtag_debug_module_translator:av_waitrequest
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata                                       : std_logic_vector(31 downto 0);  -- cpu_0_jtag_debug_module_translator:av_writedata -> cpu_0:jtag_debug_module_writedata
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address                                         : std_logic_vector(8 downto 0);   -- cpu_0_jtag_debug_module_translator:av_address -> cpu_0:jtag_debug_module_address
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write                                           : std_logic;                      -- cpu_0_jtag_debug_module_translator:av_write -> cpu_0:jtag_debug_module_write
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read                                            : std_logic;                      -- cpu_0_jtag_debug_module_translator:av_read -> cpu_0:jtag_debug_module_read
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata                                        : std_logic_vector(31 downto 0);  -- cpu_0:jtag_debug_module_readdata -> cpu_0_jtag_debug_module_translator:av_readdata
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess                                     : std_logic;                      -- cpu_0_jtag_debug_module_translator:av_debugaccess -> cpu_0:jtag_debug_module_debugaccess
	signal cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable                                      : std_logic_vector(3 downto 0);   -- cpu_0_jtag_debug_module_translator:av_byteenable -> cpu_0:jtag_debug_module_byteenable
	signal sdram_0_s1_translator_avalon_anti_slave_0_waitrequest                                                  : std_logic;                      -- sdram_0:za_waitrequest -> sdram_0_s1_translator:av_waitrequest
	signal sdram_0_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator:av_writedata -> sdram_0:az_data
	signal sdram_0_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(21 downto 0);  -- sdram_0_s1_translator:av_address -> sdram_0:az_addr
	signal sdram_0_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- sdram_0_s1_translator:av_chipselect -> sdram_0:az_cs
	signal sdram_0_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- sdram_0_s1_translator:av_write -> sdram_0_s1_translator_avalon_anti_slave_0_write:in
	signal sdram_0_s1_translator_avalon_anti_slave_0_read                                                         : std_logic;                      -- sdram_0_s1_translator:av_read -> sdram_0_s1_translator_avalon_anti_slave_0_read:in
	signal sdram_0_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(15 downto 0);  -- sdram_0:za_data -> sdram_0_s1_translator:av_readdata
	signal sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid                                                : std_logic;                      -- sdram_0:za_valid -> sdram_0_s1_translator:av_readdatavalid
	signal sdram_0_s1_translator_avalon_anti_slave_0_byteenable                                                   : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator:av_byteenable -> sdram_0_s1_translator_avalon_anti_slave_0_byteenable:in
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- epcs_controller_epcs_control_port_translator:av_writedata -> epcs_controller:writedata
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address                               : std_logic_vector(8 downto 0);   -- epcs_controller_epcs_control_port_translator:av_address -> epcs_controller:address
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect                            : std_logic;                      -- epcs_controller_epcs_control_port_translator:av_chipselect -> epcs_controller:chipselect
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- epcs_controller_epcs_control_port_translator:av_write -> epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write:in
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- epcs_controller_epcs_control_port_translator:av_read -> epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read:in
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- epcs_controller:readdata -> epcs_controller_epcs_control_port_translator:av_readdata
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest                                             : std_logic;                      -- cfi_flash_0:uas_waitrequest -> cfi_flash_0_uas_translator:av_waitrequest
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount                                              : std_logic_vector(0 downto 0);   -- cfi_flash_0_uas_translator:av_burstcount -> cfi_flash_0:uas_burstcount
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata                                               : std_logic_vector(7 downto 0);   -- cfi_flash_0_uas_translator:av_writedata -> cfi_flash_0:uas_writedata
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_address                                                 : std_logic_vector(21 downto 0);  -- cfi_flash_0_uas_translator:av_address -> cfi_flash_0:uas_address
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_lock                                                    : std_logic;                      -- cfi_flash_0_uas_translator:av_lock -> cfi_flash_0:uas_lock
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_write                                                   : std_logic;                      -- cfi_flash_0_uas_translator:av_write -> cfi_flash_0:uas_write
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_read                                                    : std_logic;                      -- cfi_flash_0_uas_translator:av_read -> cfi_flash_0:uas_read
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata                                                : std_logic_vector(7 downto 0);   -- cfi_flash_0:uas_readdata -> cfi_flash_0_uas_translator:av_readdata
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess                                             : std_logic;                      -- cfi_flash_0_uas_translator:av_debugaccess -> cfi_flash_0:uas_debugaccess
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid                                           : std_logic;                      -- cfi_flash_0:uas_readdatavalid -> cfi_flash_0_uas_translator:av_readdatavalid
	signal cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable                                              : std_logic_vector(0 downto 0);   -- cfi_flash_0_uas_translator:av_byteenable -> cfi_flash_0:uas_byteenable
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address                                      : std_logic_vector(0 downto 0);   -- sysid_qsys_0_control_slave_translator:av_address -> sysid_qsys_0:address
	signal sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata                                     : std_logic_vector(31 downto 0);  -- sysid_qsys_0:readdata -> sysid_qsys_0_control_slave_translator:av_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest                               : std_logic;                      -- jtag_uart_0:av_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator:av_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata                                 : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:av_writedata -> jtag_uart_0:av_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address                                   : std_logic_vector(0 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator:av_address -> jtag_uart_0:av_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect                                : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_chipselect -> jtag_uart_0:av_chipselect
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write                                     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_write -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read                                      : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:av_read -> jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:in
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata                                  : std_logic_vector(31 downto 0);  -- jtag_uart_0:av_readdata -> jtag_uart_0_avalon_jtag_slave_translator:av_readdata
	signal uart_0_s1_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(15 downto 0);  -- uart_0_s1_translator:av_writedata -> uart_0:writedata
	signal uart_0_s1_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(2 downto 0);   -- uart_0_s1_translator:av_address -> uart_0:address
	signal uart_0_s1_translator_avalon_anti_slave_0_chipselect                                                    : std_logic;                      -- uart_0_s1_translator:av_chipselect -> uart_0:chipselect
	signal uart_0_s1_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- uart_0_s1_translator:av_write -> uart_0_s1_translator_avalon_anti_slave_0_write:in
	signal uart_0_s1_translator_avalon_anti_slave_0_read                                                          : std_logic;                      -- uart_0_s1_translator:av_read -> uart_0_s1_translator_avalon_anti_slave_0_read:in
	signal uart_0_s1_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(15 downto 0);  -- uart_0:readdata -> uart_0_s1_translator:av_readdata
	signal uart_0_s1_translator_avalon_anti_slave_0_begintransfer                                                 : std_logic;                      -- uart_0_s1_translator:av_begintransfer -> uart_0:begintransfer
	signal timer_0_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(15 downto 0);  -- timer_0_s1_translator:av_writedata -> timer_0:writedata
	signal timer_0_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(2 downto 0);   -- timer_0_s1_translator:av_address -> timer_0:address
	signal timer_0_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- timer_0_s1_translator:av_chipselect -> timer_0:chipselect
	signal timer_0_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- timer_0_s1_translator:av_write -> timer_0_s1_translator_avalon_anti_slave_0_write:in
	signal timer_0_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(15 downto 0);  -- timer_0:readdata -> timer_0_s1_translator:av_readdata
	signal timer_1_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(15 downto 0);  -- timer_1_s1_translator:av_writedata -> timer_1:writedata
	signal timer_1_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(2 downto 0);   -- timer_1_s1_translator:av_address -> timer_1:address
	signal timer_1_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- timer_1_s1_translator:av_chipselect -> timer_1:chipselect
	signal timer_1_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- timer_1_s1_translator:av_write -> timer_1_s1_translator_avalon_anti_slave_0_write:in
	signal timer_1_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(15 downto 0);  -- timer_1:readdata -> timer_1_s1_translator:av_readdata
	signal lcd_16207_0_control_slave_translator_avalon_anti_slave_0_writedata                                     : std_logic_vector(7 downto 0);   -- lcd_16207_0_control_slave_translator:av_writedata -> lcd_16207_0:writedata
	signal lcd_16207_0_control_slave_translator_avalon_anti_slave_0_address                                       : std_logic_vector(1 downto 0);   -- lcd_16207_0_control_slave_translator:av_address -> lcd_16207_0:address
	signal lcd_16207_0_control_slave_translator_avalon_anti_slave_0_write                                         : std_logic;                      -- lcd_16207_0_control_slave_translator:av_write -> lcd_16207_0:write
	signal lcd_16207_0_control_slave_translator_avalon_anti_slave_0_read                                          : std_logic;                      -- lcd_16207_0_control_slave_translator:av_read -> lcd_16207_0:read
	signal lcd_16207_0_control_slave_translator_avalon_anti_slave_0_readdata                                      : std_logic_vector(7 downto 0);   -- lcd_16207_0:readdata -> lcd_16207_0_control_slave_translator:av_readdata
	signal lcd_16207_0_control_slave_translator_avalon_anti_slave_0_begintransfer                                 : std_logic;                      -- lcd_16207_0_control_slave_translator:av_begintransfer -> lcd_16207_0:begintransfer
	signal led_red_s1_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(31 downto 0);  -- led_red_s1_translator:av_writedata -> led_red:writedata
	signal led_red_s1_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(1 downto 0);   -- led_red_s1_translator:av_address -> led_red:address
	signal led_red_s1_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- led_red_s1_translator:av_chipselect -> led_red:chipselect
	signal led_red_s1_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- led_red_s1_translator:av_write -> led_red_s1_translator_avalon_anti_slave_0_write:in
	signal led_red_s1_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(31 downto 0);  -- led_red:readdata -> led_red_s1_translator:av_readdata
	signal led_green_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0);  -- led_green_s1_translator:av_writedata -> led_green:writedata
	signal led_green_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);   -- led_green_s1_translator:av_address -> led_green:address
	signal led_green_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                      -- led_green_s1_translator:av_chipselect -> led_green:chipselect
	signal led_green_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                      -- led_green_s1_translator:av_write -> led_green_s1_translator_avalon_anti_slave_0_write:in
	signal led_green_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0);  -- led_green:readdata -> led_green_s1_translator:av_readdata
	signal button_pio_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(31 downto 0);  -- button_pio_s1_translator:av_writedata -> button_pio:writedata
	signal button_pio_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);   -- button_pio_s1_translator:av_address -> button_pio:address
	signal button_pio_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	signal button_pio_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- button_pio_s1_translator:av_write -> button_pio_s1_translator_avalon_anti_slave_0_write:in
	signal button_pio_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- button_pio:readdata -> button_pio_s1_translator:av_readdata
	signal switch_pio_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(1 downto 0);   -- switch_pio_s1_translator:av_address -> switch_pio:address
	signal switch_pio_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(31 downto 0);  -- switch_pio:readdata -> switch_pio_s1_translator:av_readdata
	signal sd_dat_s1_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(31 downto 0);  -- SD_DAT_s1_translator:av_writedata -> SD_DAT:writedata
	signal sd_dat_s1_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(1 downto 0);   -- SD_DAT_s1_translator:av_address -> SD_DAT:address
	signal sd_dat_s1_translator_avalon_anti_slave_0_chipselect                                                    : std_logic;                      -- SD_DAT_s1_translator:av_chipselect -> SD_DAT:chipselect
	signal sd_dat_s1_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- SD_DAT_s1_translator:av_write -> sd_dat_s1_translator_avalon_anti_slave_0_write:in
	signal sd_dat_s1_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(31 downto 0);  -- SD_DAT:readdata -> SD_DAT_s1_translator:av_readdata
	signal sd_cmd_s1_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(31 downto 0);  -- SD_CMD_s1_translator:av_writedata -> SD_CMD:writedata
	signal sd_cmd_s1_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(1 downto 0);   -- SD_CMD_s1_translator:av_address -> SD_CMD:address
	signal sd_cmd_s1_translator_avalon_anti_slave_0_chipselect                                                    : std_logic;                      -- SD_CMD_s1_translator:av_chipselect -> SD_CMD:chipselect
	signal sd_cmd_s1_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- SD_CMD_s1_translator:av_write -> sd_cmd_s1_translator_avalon_anti_slave_0_write:in
	signal sd_cmd_s1_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(31 downto 0);  -- SD_CMD:readdata -> SD_CMD_s1_translator:av_readdata
	signal sd_clk_s1_translator_avalon_anti_slave_0_writedata                                                     : std_logic_vector(31 downto 0);  -- SD_CLK_s1_translator:av_writedata -> SD_CLK:writedata
	signal sd_clk_s1_translator_avalon_anti_slave_0_address                                                       : std_logic_vector(1 downto 0);   -- SD_CLK_s1_translator:av_address -> SD_CLK:address
	signal sd_clk_s1_translator_avalon_anti_slave_0_chipselect                                                    : std_logic;                      -- SD_CLK_s1_translator:av_chipselect -> SD_CLK:chipselect
	signal sd_clk_s1_translator_avalon_anti_slave_0_write                                                         : std_logic;                      -- SD_CLK_s1_translator:av_write -> sd_clk_s1_translator_avalon_anti_slave_0_write:in
	signal sd_clk_s1_translator_avalon_anti_slave_0_readdata                                                      : std_logic_vector(31 downto 0);  -- SD_CLK:readdata -> SD_CLK_s1_translator:av_readdata
	signal isp1362_hc_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(15 downto 0);  -- ISP1362_hc_translator:av_writedata -> ISP1362:avs_hc_writedata_iDATA
	signal isp1362_hc_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(0 downto 0);   -- ISP1362_hc_translator:av_address -> ISP1362:avs_hc_address_iADDR
	signal isp1362_hc_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- ISP1362_hc_translator:av_chipselect -> isp1362_hc_translator_avalon_anti_slave_0_chipselect:in
	signal isp1362_hc_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- ISP1362_hc_translator:av_write -> isp1362_hc_translator_avalon_anti_slave_0_write:in
	signal isp1362_hc_translator_avalon_anti_slave_0_read                                                         : std_logic;                      -- ISP1362_hc_translator:av_read -> isp1362_hc_translator_avalon_anti_slave_0_read:in
	signal isp1362_hc_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(15 downto 0);  -- ISP1362:avs_hc_readdata_oDATA -> ISP1362_hc_translator:av_readdata
	signal isp1362_dc_translator_avalon_anti_slave_0_writedata                                                    : std_logic_vector(15 downto 0);  -- ISP1362_dc_translator:av_writedata -> ISP1362:avs_dc_writedata_iDATA
	signal isp1362_dc_translator_avalon_anti_slave_0_address                                                      : std_logic_vector(0 downto 0);   -- ISP1362_dc_translator:av_address -> ISP1362:avs_dc_address_iADDR
	signal isp1362_dc_translator_avalon_anti_slave_0_chipselect                                                   : std_logic;                      -- ISP1362_dc_translator:av_chipselect -> isp1362_dc_translator_avalon_anti_slave_0_chipselect:in
	signal isp1362_dc_translator_avalon_anti_slave_0_write                                                        : std_logic;                      -- ISP1362_dc_translator:av_write -> isp1362_dc_translator_avalon_anti_slave_0_write:in
	signal isp1362_dc_translator_avalon_anti_slave_0_read                                                         : std_logic;                      -- ISP1362_dc_translator:av_read -> isp1362_dc_translator_avalon_anti_slave_0_read:in
	signal isp1362_dc_translator_avalon_anti_slave_0_readdata                                                     : std_logic_vector(15 downto 0);  -- ISP1362:avs_dc_readdata_oDATA -> ISP1362_dc_translator:av_readdata
	signal audio_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(15 downto 0);  -- Audio_0_avalon_slave_0_translator:av_writedata -> Audio_0:iDATA
	signal audio_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                            : std_logic;                      -- Audio_0_avalon_slave_0_translator:av_write -> Audio_0:iWR
	signal audio_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(15 downto 0);  -- Audio_0:oDATA -> Audio_0_avalon_slave_0_translator:av_readdata
	signal vga_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                          : std_logic_vector(15 downto 0);  -- VGA_0_avalon_slave_0_translator:av_writedata -> VGA_0:iDATA
	signal vga_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                            : std_logic_vector(18 downto 0);  -- VGA_0_avalon_slave_0_translator:av_address -> VGA_0:iADDR
	signal vga_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                                         : std_logic;                      -- VGA_0_avalon_slave_0_translator:av_chipselect -> VGA_0:iCS
	signal vga_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                              : std_logic;                      -- VGA_0_avalon_slave_0_translator:av_write -> VGA_0:iWR
	signal vga_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                               : std_logic;                      -- VGA_0_avalon_slave_0_translator:av_read -> VGA_0:iRD
	signal vga_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                           : std_logic_vector(15 downto 0);  -- VGA_0:oDATA -> VGA_0_avalon_slave_0_translator:av_readdata
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                        : std_logic_vector(15 downto 0);  -- DM9000A_avalon_slave_0_translator:av_writedata -> DM9000A:iDATA
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address                                          : std_logic_vector(0 downto 0);   -- DM9000A_avalon_slave_0_translator:av_address -> DM9000A:iCMD
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                                       : std_logic;                      -- DM9000A_avalon_slave_0_translator:av_chipselect -> dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect:in
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write                                            : std_logic;                      -- DM9000A_avalon_slave_0_translator:av_write -> dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write:in
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read                                             : std_logic;                      -- DM9000A_avalon_slave_0_translator:av_read -> dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read:in
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                         : std_logic_vector(15 downto 0);  -- DM9000A:oDATA -> DM9000A_avalon_slave_0_translator:av_readdata
	signal seg7_display_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0);  -- SEG7_Display_avalon_slave_0_translator:av_writedata -> SEG7_Display:iDIG
	signal seg7_display_avalon_slave_0_translator_avalon_anti_slave_0_write                                       : std_logic;                      -- SEG7_Display_avalon_slave_0_translator:av_write -> SEG7_Display:iWR
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                         : std_logic_vector(15 downto 0);  -- sram_0_avalon_slave_0_translator:av_writedata -> sram_0:iDATA
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                           : std_logic_vector(17 downto 0);  -- sram_0_avalon_slave_0_translator:av_address -> sram_0:iADDR
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                                        : std_logic;                      -- sram_0_avalon_slave_0_translator:av_chipselect -> sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect:in
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                             : std_logic;                      -- sram_0_avalon_slave_0_translator:av_write -> sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write:in
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                              : std_logic;                      -- sram_0_avalon_slave_0_translator:av_read -> sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read:in
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                          : std_logic_vector(15 downto 0);  -- sram_0:oDATA -> sram_0_avalon_slave_0_translator:av_readdata
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable                                        : std_logic_vector(1 downto 0);   -- sram_0_avalon_slave_0_translator:av_byteenable -> sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable:in
	signal lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                                   : std_logic_vector(31 downto 0);  -- lab7_FINAL_0_avalon_slave_0_translator:av_writedata -> lab7_FINAL_0:writedata
	signal lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_address                                     : std_logic_vector(0 downto 0);   -- lab7_FINAL_0_avalon_slave_0_translator:av_address -> lab7_FINAL_0:add
	signal lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                                  : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator:av_chipselect -> lab7_FINAL_0:chipselect
	signal lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                       : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator:av_write -> lab7_FINAL_0:write_en
	signal lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                        : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator:av_read -> lab7_FINAL_0:read_en
	signal lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                                    : std_logic_vector(31 downto 0);  -- lab7_FINAL_0:readdata -> lab7_FINAL_0_avalon_slave_0_translator:av_readdata
	signal motor_cw_s1_translator_avalon_anti_slave_0_writedata                                                   : std_logic_vector(31 downto 0);  -- motor_cw_s1_translator:av_writedata -> motor_cw:writedata
	signal motor_cw_s1_translator_avalon_anti_slave_0_address                                                     : std_logic_vector(1 downto 0);   -- motor_cw_s1_translator:av_address -> motor_cw:address
	signal motor_cw_s1_translator_avalon_anti_slave_0_chipselect                                                  : std_logic;                      -- motor_cw_s1_translator:av_chipselect -> motor_cw:chipselect
	signal motor_cw_s1_translator_avalon_anti_slave_0_write                                                       : std_logic;                      -- motor_cw_s1_translator:av_write -> motor_cw_s1_translator_avalon_anti_slave_0_write:in
	signal motor_cw_s1_translator_avalon_anti_slave_0_readdata                                                    : std_logic_vector(31 downto 0);  -- motor_cw:readdata -> motor_cw_s1_translator:av_readdata
	signal motor_ccw_s1_translator_avalon_anti_slave_0_writedata                                                  : std_logic_vector(31 downto 0);  -- motor_ccw_s1_translator:av_writedata -> motor_ccw:writedata
	signal motor_ccw_s1_translator_avalon_anti_slave_0_address                                                    : std_logic_vector(1 downto 0);   -- motor_ccw_s1_translator:av_address -> motor_ccw:address
	signal motor_ccw_s1_translator_avalon_anti_slave_0_chipselect                                                 : std_logic;                      -- motor_ccw_s1_translator:av_chipselect -> motor_ccw:chipselect
	signal motor_ccw_s1_translator_avalon_anti_slave_0_write                                                      : std_logic;                      -- motor_ccw_s1_translator:av_write -> motor_ccw_s1_translator_avalon_anti_slave_0_write:in
	signal motor_ccw_s1_translator_avalon_anti_slave_0_readdata                                                   : std_logic_vector(31 downto 0);  -- motor_ccw:readdata -> motor_ccw_s1_translator:av_readdata
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest                              : std_logic;                      -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_instruction_master_translator:uav_waitrequest
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount                               : std_logic_vector(2 downto 0);   -- cpu_0_instruction_master_translator:uav_burstcount -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_writedata                                : std_logic_vector(31 downto 0);  -- cpu_0_instruction_master_translator:uav_writedata -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_address                                  : std_logic_vector(24 downto 0);  -- cpu_0_instruction_master_translator:uav_address -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_lock                                     : std_logic;                      -- cpu_0_instruction_master_translator:uav_lock -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_write                                    : std_logic;                      -- cpu_0_instruction_master_translator:uav_write -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_read                                     : std_logic;                      -- cpu_0_instruction_master_translator:uav_read -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_readdata                                 : std_logic_vector(31 downto 0);  -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_instruction_master_translator:uav_readdata
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess                              : std_logic;                      -- cpu_0_instruction_master_translator:uav_debugaccess -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable                               : std_logic_vector(3 downto 0);   -- cpu_0_instruction_master_translator:uav_byteenable -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid                            : std_logic;                      -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_instruction_master_translator:uav_readdatavalid
	signal cpu_0_data_master_translator_avalon_universal_master_0_waitrequest                                     : std_logic;                      -- cpu_0_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_0_data_master_translator:uav_waitrequest
	signal cpu_0_data_master_translator_avalon_universal_master_0_burstcount                                      : std_logic_vector(2 downto 0);   -- cpu_0_data_master_translator:uav_burstcount -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_0_data_master_translator_avalon_universal_master_0_writedata                                       : std_logic_vector(31 downto 0);  -- cpu_0_data_master_translator:uav_writedata -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_0_data_master_translator_avalon_universal_master_0_address                                         : std_logic_vector(24 downto 0);  -- cpu_0_data_master_translator:uav_address -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_0_data_master_translator_avalon_universal_master_0_lock                                            : std_logic;                      -- cpu_0_data_master_translator:uav_lock -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_0_data_master_translator_avalon_universal_master_0_write                                           : std_logic;                      -- cpu_0_data_master_translator:uav_write -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_0_data_master_translator_avalon_universal_master_0_read                                            : std_logic;                      -- cpu_0_data_master_translator:uav_read -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_0_data_master_translator_avalon_universal_master_0_readdata                                        : std_logic_vector(31 downto 0);  -- cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_0_data_master_translator:uav_readdata
	signal cpu_0_data_master_translator_avalon_universal_master_0_debugaccess                                     : std_logic;                      -- cpu_0_data_master_translator:uav_debugaccess -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_0_data_master_translator_avalon_universal_master_0_byteenable                                      : std_logic_vector(3 downto 0);   -- cpu_0_data_master_translator:uav_byteenable -> cpu_0_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid                                   : std_logic;                      -- cpu_0_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_0_data_master_translator:uav_readdatavalid
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest                       : std_logic;                      -- cpu_0_jtag_debug_module_translator:uav_waitrequest -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount                        : std_logic_vector(2 downto 0);   -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_burstcount -> cpu_0_jtag_debug_module_translator:uav_burstcount
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata                         : std_logic_vector(31 downto 0);  -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_writedata -> cpu_0_jtag_debug_module_translator:uav_writedata
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address                           : std_logic_vector(24 downto 0);  -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_address -> cpu_0_jtag_debug_module_translator:uav_address
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write                             : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_write -> cpu_0_jtag_debug_module_translator:uav_write
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock                              : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_lock -> cpu_0_jtag_debug_module_translator:uav_lock
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read                              : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_read -> cpu_0_jtag_debug_module_translator:uav_read
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata                          : std_logic_vector(31 downto 0);  -- cpu_0_jtag_debug_module_translator:uav_readdata -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid                     : std_logic;                      -- cpu_0_jtag_debug_module_translator:uav_readdatavalid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess                       : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cpu_0_jtag_debug_module_translator:uav_debugaccess
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable                        : std_logic_vector(3 downto 0);   -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:m0_byteenable -> cpu_0_jtag_debug_module_translator:uav_byteenable
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid                      : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket              : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data                       : std_logic_vector(102 downto 0); -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready                      : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket             : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                   : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket           : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                    : std_logic_vector(102 downto 0); -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                   : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                 : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                  : std_logic_vector(33 downto 0);  -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                 : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- sdram_0_s1_translator:uav_waitrequest -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_0_s1_translator:uav_burstcount
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_0_s1_translator:uav_writedata
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_0_s1_translator:uav_address
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_0_s1_translator:uav_write
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_0_s1_translator:uav_lock
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_0_s1_translator:uav_read
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(15 downto 0);  -- sdram_0_s1_translator:uav_readdata -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- sdram_0_s1_translator:uav_readdatavalid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_0_s1_translator:uav_debugaccess
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_0_s1_translator:uav_byteenable
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(84 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(84 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(17 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                              : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                               : std_logic_vector(17 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                              : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- epcs_controller_epcs_control_port_translator:uav_waitrequest -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_burstcount -> epcs_controller_epcs_control_port_translator:uav_burstcount
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_writedata -> epcs_controller_epcs_control_port_translator:uav_writedata
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(24 downto 0);  -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_address -> epcs_controller_epcs_control_port_translator:uav_address
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_write -> epcs_controller_epcs_control_port_translator:uav_write
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_lock -> epcs_controller_epcs_control_port_translator:uav_lock
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_read -> epcs_controller_epcs_control_port_translator:uav_read
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- epcs_controller_epcs_control_port_translator:uav_readdata -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdata
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- epcs_controller_epcs_control_port_translator:uav_readdatavalid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_debugaccess -> epcs_controller_epcs_control_port_translator:uav_debugaccess
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:m0_byteenable -> epcs_controller_epcs_control_port_translator:uav_byteenable
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(102 downto 0); -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(102 downto 0); -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rf_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest                               : std_logic;                      -- cfi_flash_0_uas_translator:uav_waitrequest -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount                                : std_logic_vector(0 downto 0);   -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_burstcount -> cfi_flash_0_uas_translator:uav_burstcount
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata                                 : std_logic_vector(7 downto 0);   -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_writedata -> cfi_flash_0_uas_translator:uav_writedata
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address                                   : std_logic_vector(24 downto 0);  -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_address -> cfi_flash_0_uas_translator:uav_address
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write                                     : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_write -> cfi_flash_0_uas_translator:uav_write
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock                                      : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_lock -> cfi_flash_0_uas_translator:uav_lock
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read                                      : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_read -> cfi_flash_0_uas_translator:uav_read
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata                                  : std_logic_vector(7 downto 0);   -- cfi_flash_0_uas_translator:uav_readdata -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdata
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid                             : std_logic;                      -- cfi_flash_0_uas_translator:uav_readdatavalid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess                               : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_debugaccess -> cfi_flash_0_uas_translator:uav_debugaccess
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable                                : std_logic_vector(0 downto 0);   -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:m0_byteenable -> cfi_flash_0_uas_translator:uav_byteenable
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                        : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid                              : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                      : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data                               : std_logic_vector(75 downto 0);  -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready                              : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                     : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                           : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                   : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                            : std_logic_vector(75 downto 0);  -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                           : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rf_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                         : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                          : std_logic_vector(9 downto 0);   -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                         : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid                         : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data                          : std_logic_vector(9 downto 0);   -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready                         : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                    : std_logic;                      -- sysid_qsys_0_control_slave_translator:uav_waitrequest -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                     : std_logic_vector(2 downto 0);   -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> sysid_qsys_0_control_slave_translator:uav_burstcount
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                      : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> sysid_qsys_0_control_slave_translator:uav_writedata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address                        : std_logic_vector(24 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> sysid_qsys_0_control_slave_translator:uav_address
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write                          : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> sysid_qsys_0_control_slave_translator:uav_write
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                           : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> sysid_qsys_0_control_slave_translator:uav_lock
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read                           : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> sysid_qsys_0_control_slave_translator:uav_read
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                       : std_logic_vector(31 downto 0);  -- sysid_qsys_0_control_slave_translator:uav_readdata -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                  : std_logic;                      -- sysid_qsys_0_control_slave_translator:uav_readdatavalid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                    : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sysid_qsys_0_control_slave_translator:uav_debugaccess
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                     : std_logic_vector(3 downto 0);   -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> sysid_qsys_0_control_slave_translator:uav_byteenable
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket             : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                   : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket           : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                    : std_logic_vector(102 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                   : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket          : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket        : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                 : std_logic_vector(102 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid              : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data               : std_logic_vector(33 downto 0);  -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready              : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                  : std_logic_vector(2 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_0_avalon_jtag_slave_translator:uav_burstcount
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata                   : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_0_avalon_jtag_slave_translator:uav_writedata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address                     : std_logic_vector(24 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_0_avalon_jtag_slave_translator:uav_address
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_0_avalon_jtag_slave_translator:uav_write
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_0_avalon_jtag_slave_translator:uav_lock
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read                        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_0_avalon_jtag_slave_translator:uav_read
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata                    : std_logic_vector(31 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_0_avalon_jtag_slave_translator:uav_debugaccess
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                  : std_logic_vector(3 downto 0);   -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_0_avalon_jtag_slave_translator:uav_byteenable
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket          : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket        : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data                 : std_logic_vector(102 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid             : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket     : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data              : std_logic_vector(102 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready             : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data            : std_logic_vector(33 downto 0);  -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- uart_0_s1_translator:uav_waitrequest -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> uart_0_s1_translator:uav_burstcount
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> uart_0_s1_translator:uav_writedata
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(24 downto 0);  -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> uart_0_s1_translator:uav_address
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> uart_0_s1_translator:uav_write
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> uart_0_s1_translator:uav_lock
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> uart_0_s1_translator:uav_read
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- uart_0_s1_translator:uav_readdata -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- uart_0_s1_translator:uav_readdatavalid -> uart_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> uart_0_s1_translator:uav_debugaccess
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- uart_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> uart_0_s1_translator:uav_byteenable
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(102 downto 0); -- uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(102 downto 0); -- uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(33 downto 0);  -- uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- timer_0_s1_translator:uav_waitrequest -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_0_s1_translator:uav_burstcount
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_0_s1_translator:uav_writedata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_0_s1_translator:uav_address
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_0_s1_translator:uav_write
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_0_s1_translator:uav_lock
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_0_s1_translator:uav_read
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- timer_0_s1_translator:uav_readdata -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- timer_0_s1_translator:uav_readdatavalid -> timer_0_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_0_s1_translator:uav_debugaccess
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- timer_0_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_0_s1_translator:uav_byteenable
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(102 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(102 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- timer_1_s1_translator:uav_waitrequest -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> timer_1_s1_translator:uav_burstcount
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> timer_1_s1_translator:uav_writedata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_address -> timer_1_s1_translator:uav_address
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_write -> timer_1_s1_translator:uav_write
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_lock -> timer_1_s1_translator:uav_lock
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_read -> timer_1_s1_translator:uav_read
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- timer_1_s1_translator:uav_readdata -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- timer_1_s1_translator:uav_readdatavalid -> timer_1_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> timer_1_s1_translator:uav_debugaccess
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- timer_1_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> timer_1_s1_translator:uav_byteenable
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(102 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(102 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest                     : std_logic;                      -- lcd_16207_0_control_slave_translator:uav_waitrequest -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount                      : std_logic_vector(2 downto 0);   -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> lcd_16207_0_control_slave_translator:uav_burstcount
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata                       : std_logic_vector(31 downto 0);  -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> lcd_16207_0_control_slave_translator:uav_writedata
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address                         : std_logic_vector(24 downto 0);  -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_address -> lcd_16207_0_control_slave_translator:uav_address
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write                           : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_write -> lcd_16207_0_control_slave_translator:uav_write
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock                            : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_lock -> lcd_16207_0_control_slave_translator:uav_lock
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read                            : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_read -> lcd_16207_0_control_slave_translator:uav_read
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata                        : std_logic_vector(31 downto 0);  -- lcd_16207_0_control_slave_translator:uav_readdata -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid                   : std_logic;                      -- lcd_16207_0_control_slave_translator:uav_readdatavalid -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess                     : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lcd_16207_0_control_slave_translator:uav_debugaccess
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable                      : std_logic_vector(3 downto 0);   -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> lcd_16207_0_control_slave_translator:uav_byteenable
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket              : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid                    : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket            : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data                     : std_logic_vector(102 downto 0); -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready                    : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket           : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                 : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket         : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                  : std_logic_vector(102 downto 0); -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                 : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid               : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                : std_logic_vector(33 downto 0);  -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready               : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- led_red_s1_translator:uav_waitrequest -> led_red_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_red_s1_translator:uav_burstcount
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_red_s1_translator:uav_writedata
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_red_s1_translator:uav_address
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_red_s1_translator:uav_write
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_red_s1_translator:uav_lock
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_red_s1_translator:uav_read
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- led_red_s1_translator:uav_readdata -> led_red_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- led_red_s1_translator:uav_readdatavalid -> led_red_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_red_s1_translator:uav_debugaccess
	signal led_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- led_red_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_red_s1_translator:uav_byteenable
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(102 downto 0); -- led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(102 downto 0); -- led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_red_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- led_green_s1_translator:uav_waitrequest -> led_green_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);   -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_green_s1_translator:uav_burstcount
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0);  -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_green_s1_translator:uav_writedata
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(24 downto 0);  -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_green_s1_translator:uav_address
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_green_s1_translator:uav_write
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_green_s1_translator:uav_lock
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_green_s1_translator:uav_read
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0);  -- led_green_s1_translator:uav_readdata -> led_green_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- led_green_s1_translator:uav_readdatavalid -> led_green_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_green_s1_translator:uav_debugaccess
	signal led_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);   -- led_green_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_green_s1_translator:uav_byteenable
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(102 downto 0); -- led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(102 downto 0); -- led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0);  -- led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_green_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(24 downto 0);  -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(102 downto 0); -- button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(102 downto 0); -- button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- switch_pio_s1_translator:uav_waitrequest -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(2 downto 0);   -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> switch_pio_s1_translator:uav_burstcount
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(31 downto 0);  -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> switch_pio_s1_translator:uav_writedata
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(24 downto 0);  -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> switch_pio_s1_translator:uav_address
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> switch_pio_s1_translator:uav_write
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> switch_pio_s1_translator:uav_lock
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> switch_pio_s1_translator:uav_read
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(31 downto 0);  -- switch_pio_s1_translator:uav_readdata -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- switch_pio_s1_translator:uav_readdatavalid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> switch_pio_s1_translator:uav_debugaccess
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(3 downto 0);   -- switch_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> switch_pio_s1_translator:uav_byteenable
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(102 downto 0); -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(102 downto 0); -- switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(33 downto 0);  -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- SD_DAT_s1_translator:uav_waitrequest -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_DAT_s1_translator:uav_burstcount
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_DAT_s1_translator:uav_writedata
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(24 downto 0);  -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_DAT_s1_translator:uav_address
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_DAT_s1_translator:uav_write
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_DAT_s1_translator:uav_lock
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_DAT_s1_translator:uav_read
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- SD_DAT_s1_translator:uav_readdata -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- SD_DAT_s1_translator:uav_readdatavalid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_DAT_s1_translator:uav_debugaccess
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_DAT_s1_translator:uav_byteenable
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(102 downto 0); -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(102 downto 0); -- SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(33 downto 0);  -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- SD_CMD_s1_translator:uav_waitrequest -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_CMD_s1_translator:uav_burstcount
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_CMD_s1_translator:uav_writedata
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(24 downto 0);  -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_CMD_s1_translator:uav_address
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_CMD_s1_translator:uav_write
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_CMD_s1_translator:uav_lock
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_CMD_s1_translator:uav_read
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- SD_CMD_s1_translator:uav_readdata -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- SD_CMD_s1_translator:uav_readdatavalid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_CMD_s1_translator:uav_debugaccess
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_CMD_s1_translator:uav_byteenable
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(102 downto 0); -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(102 downto 0); -- SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(33 downto 0);  -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                     : std_logic;                      -- SD_CLK_s1_translator:uav_waitrequest -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                      : std_logic_vector(2 downto 0);   -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> SD_CLK_s1_translator:uav_burstcount
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                       : std_logic_vector(31 downto 0);  -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> SD_CLK_s1_translator:uav_writedata
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address                                         : std_logic_vector(24 downto 0);  -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_address -> SD_CLK_s1_translator:uav_address
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write                                           : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_write -> SD_CLK_s1_translator:uav_write
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock                                            : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_lock -> SD_CLK_s1_translator:uav_lock
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read                                            : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_read -> SD_CLK_s1_translator:uav_read
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                        : std_logic_vector(31 downto 0);  -- SD_CLK_s1_translator:uav_readdata -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                   : std_logic;                      -- SD_CLK_s1_translator:uav_readdatavalid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                     : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SD_CLK_s1_translator:uav_debugaccess
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                      : std_logic_vector(3 downto 0);   -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> SD_CLK_s1_translator:uav_byteenable
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                              : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                    : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                            : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                     : std_logic_vector(102 downto 0); -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                    : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                           : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                 : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                         : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                  : std_logic_vector(102 downto 0); -- SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                 : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                               : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                                : std_logic_vector(33 downto 0);  -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                               : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- ISP1362_hc_translator:uav_waitrequest -> ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1362_hc_translator:uav_burstcount
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1362_hc_translator:uav_writedata
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_address -> ISP1362_hc_translator:uav_address
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_write -> ISP1362_hc_translator:uav_write
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1362_hc_translator:uav_lock
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_read -> ISP1362_hc_translator:uav_read
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- ISP1362_hc_translator:uav_readdata -> ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_readdata
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- ISP1362_hc_translator:uav_readdatavalid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1362_hc_translator:uav_debugaccess
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- ISP1362_hc_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1362_hc_translator:uav_byteenable
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(102 downto 0); -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(102 downto 0); -- ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest                                    : std_logic;                      -- ISP1362_dc_translator:uav_waitrequest -> ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_burstcount                                     : std_logic_vector(2 downto 0);   -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_burstcount -> ISP1362_dc_translator:uav_burstcount
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_writedata                                      : std_logic_vector(31 downto 0);  -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_writedata -> ISP1362_dc_translator:uav_writedata
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_address                                        : std_logic_vector(24 downto 0);  -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_address -> ISP1362_dc_translator:uav_address
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_write                                          : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_write -> ISP1362_dc_translator:uav_write
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_lock                                           : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_lock -> ISP1362_dc_translator:uav_lock
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_read                                           : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_read -> ISP1362_dc_translator:uav_read
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdata                                       : std_logic_vector(31 downto 0);  -- ISP1362_dc_translator:uav_readdata -> ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_readdata
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                  : std_logic;                      -- ISP1362_dc_translator:uav_readdatavalid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess                                    : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_debugaccess -> ISP1362_dc_translator:uav_debugaccess
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_m0_byteenable                                     : std_logic_vector(3 downto 0);   -- ISP1362_dc_translator_avalon_universal_slave_0_agent:m0_byteenable -> ISP1362_dc_translator:uav_byteenable
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                             : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_valid                                   : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                           : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_data                                    : std_logic_vector(102 downto 0); -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_ready                                   : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                          : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                                : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                        : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                 : std_logic_vector(102 downto 0); -- ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                                : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rf_sink_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                              : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                               : std_logic_vector(33 downto 0);  -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                              : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- Audio_0_avalon_slave_0_translator:uav_waitrequest -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> Audio_0_avalon_slave_0_translator:uav_burstcount
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> Audio_0_avalon_slave_0_translator:uav_writedata
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(24 downto 0);  -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> Audio_0_avalon_slave_0_translator:uav_address
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> Audio_0_avalon_slave_0_translator:uav_write
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> Audio_0_avalon_slave_0_translator:uav_lock
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> Audio_0_avalon_slave_0_translator:uav_read
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- Audio_0_avalon_slave_0_translator:uav_readdata -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- Audio_0_avalon_slave_0_translator:uav_readdatavalid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> Audio_0_avalon_slave_0_translator:uav_debugaccess
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> Audio_0_avalon_slave_0_translator:uav_byteenable
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(102 downto 0); -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(102 downto 0); -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                          : std_logic;                      -- VGA_0_avalon_slave_0_translator:uav_waitrequest -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                           : std_logic_vector(2 downto 0);   -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> VGA_0_avalon_slave_0_translator:uav_burstcount
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                            : std_logic_vector(31 downto 0);  -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> VGA_0_avalon_slave_0_translator:uav_writedata
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                              : std_logic_vector(24 downto 0);  -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> VGA_0_avalon_slave_0_translator:uav_address
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                                : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> VGA_0_avalon_slave_0_translator:uav_write
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                                 : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> VGA_0_avalon_slave_0_translator:uav_lock
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                                 : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> VGA_0_avalon_slave_0_translator:uav_read
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                             : std_logic_vector(31 downto 0);  -- VGA_0_avalon_slave_0_translator:uav_readdata -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                        : std_logic;                      -- VGA_0_avalon_slave_0_translator:uav_readdatavalid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                          : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> VGA_0_avalon_slave_0_translator:uav_debugaccess
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                           : std_logic_vector(3 downto 0);   -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> VGA_0_avalon_slave_0_translator:uav_byteenable
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                   : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                         : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                 : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                          : std_logic_vector(102 downto 0); -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                         : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                      : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket              : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                       : std_logic_vector(102 downto 0); -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                      : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                    : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                     : std_logic_vector(33 downto 0);  -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                    : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                        : std_logic;                      -- DM9000A_avalon_slave_0_translator:uav_waitrequest -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                         : std_logic_vector(2 downto 0);   -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> DM9000A_avalon_slave_0_translator:uav_burstcount
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                          : std_logic_vector(31 downto 0);  -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> DM9000A_avalon_slave_0_translator:uav_writedata
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                            : std_logic_vector(24 downto 0);  -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> DM9000A_avalon_slave_0_translator:uav_address
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                              : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> DM9000A_avalon_slave_0_translator:uav_write
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                               : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> DM9000A_avalon_slave_0_translator:uav_lock
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                               : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> DM9000A_avalon_slave_0_translator:uav_read
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                           : std_logic_vector(31 downto 0);  -- DM9000A_avalon_slave_0_translator:uav_readdata -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                      : std_logic;                      -- DM9000A_avalon_slave_0_translator:uav_readdatavalid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                        : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> DM9000A_avalon_slave_0_translator:uav_debugaccess
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                         : std_logic_vector(3 downto 0);   -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> DM9000A_avalon_slave_0_translator:uav_byteenable
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                 : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                       : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket               : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                        : std_logic_vector(102 downto 0); -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                       : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket              : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                    : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket            : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                     : std_logic_vector(102 downto 0); -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                    : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                  : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                   : std_logic_vector(33 downto 0);  -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                  : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                      -- SEG7_Display_avalon_slave_0_translator:uav_waitrequest -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);   -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> SEG7_Display_avalon_slave_0_translator:uav_burstcount
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0);  -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> SEG7_Display_avalon_slave_0_translator:uav_writedata
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(24 downto 0);  -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> SEG7_Display_avalon_slave_0_translator:uav_address
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> SEG7_Display_avalon_slave_0_translator:uav_write
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> SEG7_Display_avalon_slave_0_translator:uav_lock
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> SEG7_Display_avalon_slave_0_translator:uav_read
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0);  -- SEG7_Display_avalon_slave_0_translator:uav_readdata -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                      -- SEG7_Display_avalon_slave_0_translator:uav_readdatavalid -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> SEG7_Display_avalon_slave_0_translator:uav_debugaccess
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);   -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> SEG7_Display_avalon_slave_0_translator:uav_byteenable
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(102 downto 0); -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(102 downto 0); -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0);  -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                         : std_logic;                      -- sram_0_avalon_slave_0_translator:uav_waitrequest -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                          : std_logic_vector(1 downto 0);   -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> sram_0_avalon_slave_0_translator:uav_burstcount
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                           : std_logic_vector(15 downto 0);  -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> sram_0_avalon_slave_0_translator:uav_writedata
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                             : std_logic_vector(24 downto 0);  -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> sram_0_avalon_slave_0_translator:uav_address
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                               : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> sram_0_avalon_slave_0_translator:uav_write
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                                : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> sram_0_avalon_slave_0_translator:uav_lock
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                                : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> sram_0_avalon_slave_0_translator:uav_read
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                            : std_logic_vector(15 downto 0);  -- sram_0_avalon_slave_0_translator:uav_readdata -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                       : std_logic;                      -- sram_0_avalon_slave_0_translator:uav_readdatavalid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                         : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sram_0_avalon_slave_0_translator:uav_debugaccess
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                          : std_logic_vector(1 downto 0);   -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> sram_0_avalon_slave_0_translator:uav_byteenable
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                  : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                        : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                         : std_logic_vector(84 downto 0);  -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                        : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket               : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                     : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket             : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                      : std_logic_vector(84 downto 0);  -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                     : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                   : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                    : std_logic_vector(17 downto 0);  -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                   : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest                   : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator:uav_waitrequest -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount                    : std_logic_vector(2 downto 0);   -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> lab7_FINAL_0_avalon_slave_0_translator:uav_burstcount
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata                     : std_logic_vector(31 downto 0);  -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> lab7_FINAL_0_avalon_slave_0_translator:uav_writedata
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                       : std_logic_vector(24 downto 0);  -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> lab7_FINAL_0_avalon_slave_0_translator:uav_address
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                         : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> lab7_FINAL_0_avalon_slave_0_translator:uav_write
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                          : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> lab7_FINAL_0_avalon_slave_0_translator:uav_lock
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                          : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> lab7_FINAL_0_avalon_slave_0_translator:uav_read
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                      : std_logic_vector(31 downto 0);  -- lab7_FINAL_0_avalon_slave_0_translator:uav_readdata -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid                 : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator:uav_readdatavalid -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess                   : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> lab7_FINAL_0_avalon_slave_0_translator:uav_debugaccess
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable                    : std_logic_vector(3 downto 0);   -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> lab7_FINAL_0_avalon_slave_0_translator:uav_byteenable
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket            : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid                  : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket          : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data                   : std_logic_vector(102 downto 0); -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready                  : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket         : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid               : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket       : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                : std_logic_vector(102 downto 0); -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready               : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid             : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data              : std_logic_vector(33 downto 0);  -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready             : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                   : std_logic;                      -- motor_cw_s1_translator:uav_waitrequest -> motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                    : std_logic_vector(2 downto 0);   -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> motor_cw_s1_translator:uav_burstcount
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                     : std_logic_vector(31 downto 0);  -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> motor_cw_s1_translator:uav_writedata
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_address                                       : std_logic_vector(24 downto 0);  -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_address -> motor_cw_s1_translator:uav_address
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_write                                         : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_write -> motor_cw_s1_translator:uav_write
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_lock                                          : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> motor_cw_s1_translator:uav_lock
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_read                                          : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_read -> motor_cw_s1_translator:uav_read
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                      : std_logic_vector(31 downto 0);  -- motor_cw_s1_translator:uav_readdata -> motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                 : std_logic;                      -- motor_cw_s1_translator:uav_readdatavalid -> motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                   : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> motor_cw_s1_translator:uav_debugaccess
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                    : std_logic_vector(3 downto 0);   -- motor_cw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> motor_cw_s1_translator:uav_byteenable
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                            : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                  : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                          : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                   : std_logic_vector(102 downto 0); -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                  : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                         : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                               : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                       : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                                : std_logic_vector(102 downto 0); -- motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                               : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                             : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                              : std_logic_vector(33 downto 0);  -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                             : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                  : std_logic;                      -- motor_ccw_s1_translator:uav_waitrequest -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                   : std_logic_vector(2 downto 0);   -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> motor_ccw_s1_translator:uav_burstcount
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                    : std_logic_vector(31 downto 0);  -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> motor_ccw_s1_translator:uav_writedata
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_address                                      : std_logic_vector(24 downto 0);  -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_address -> motor_ccw_s1_translator:uav_address
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_write                                        : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_write -> motor_ccw_s1_translator:uav_write
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_lock                                         : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_lock -> motor_ccw_s1_translator:uav_lock
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_read                                         : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_read -> motor_ccw_s1_translator:uav_read
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                     : std_logic_vector(31 downto 0);  -- motor_ccw_s1_translator:uav_readdata -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                                : std_logic;                      -- motor_ccw_s1_translator:uav_readdatavalid -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                  : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> motor_ccw_s1_translator:uav_debugaccess
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                   : std_logic_vector(3 downto 0);   -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> motor_ccw_s1_translator:uav_byteenable
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                           : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                 : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                         : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                  : std_logic_vector(102 downto 0); -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                 : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                        : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                              : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                      : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                               : std_logic_vector(102 downto 0); -- motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                              : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                            : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                             : std_logic_vector(33 downto 0);  -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                            : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                     : std_logic;                      -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                           : std_logic;                      -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                   : std_logic;                      -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data                            : std_logic_vector(101 downto 0); -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                           : std_logic;                      -- addr_router:sink_ready -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                            : std_logic;                      -- cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid                                  : std_logic;                      -- cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                          : std_logic;                      -- cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data                                   : std_logic_vector(101 downto 0); -- cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready                                  : std_logic;                      -- addr_router_001:sink_ready -> cpu_0_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket                       : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid                             : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket                     : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data                              : std_logic_vector(101 downto 0); -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready                             : std_logic;                      -- id_router:sink_ready -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:rp_ready
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(83 downto 0);  -- sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_001:sink_ready -> sdram_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(101 downto 0); -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	signal epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_002:sink_ready -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:rp_ready
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket                               : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid                                     : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket                             : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data                                      : std_logic_vector(74 downto 0);  -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	signal cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready                                     : std_logic;                      -- id_router_003:sink_ready -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:rp_ready
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                    : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                          : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                  : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data                           : std_logic_vector(101 downto 0); -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	signal sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                          : std_logic;                      -- id_router_004:sink_ready -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                 : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid                       : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket               : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data                        : std_logic_vector(101 downto 0); -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready                       : std_logic;                      -- id_router_005:sink_ready -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(101 downto 0); -- uart_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	signal uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_006:sink_ready -> uart_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(101 downto 0); -- timer_0_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	signal timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_007:sink_ready -> timer_0_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(101 downto 0); -- timer_1_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	signal timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_008:sink_ready -> timer_1_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket                     : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid                           : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket                   : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data                            : std_logic_vector(101 downto 0); -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	signal lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready                           : std_logic;                      -- id_router_009:sink_ready -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:rp_ready
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(101 downto 0); -- led_red_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	signal led_red_s1_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_010:sink_ready -> led_red_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_011:sink_endofpacket
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_011:sink_valid
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_011:sink_startofpacket
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(101 downto 0); -- led_green_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_011:sink_data
	signal led_green_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_011:sink_ready -> led_green_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_012:sink_endofpacket
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_012:sink_valid
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_012:sink_startofpacket
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(101 downto 0); -- button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_012:sink_data
	signal button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_012:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_013:sink_endofpacket
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_013:sink_valid
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_013:sink_startofpacket
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(101 downto 0); -- switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_013:sink_data
	signal switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router_013:sink_ready -> switch_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_014:sink_endofpacket
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_014:sink_valid
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_014:sink_startofpacket
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(101 downto 0); -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_014:sink_data
	signal sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_014:sink_ready -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_015:sink_endofpacket
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_015:sink_valid
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_015:sink_startofpacket
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(101 downto 0); -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_015:sink_data
	signal sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_015:sink_ready -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                     : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_016:sink_endofpacket
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid                                           : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_016:sink_valid
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                   : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_016:sink_startofpacket
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data                                            : std_logic_vector(101 downto 0); -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_016:sink_data
	signal sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready                                           : std_logic;                      -- id_router_016:sink_ready -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_017:sink_endofpacket
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_017:sink_valid
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_017:sink_startofpacket
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(101 downto 0); -- ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_data -> id_router_017:sink_data
	signal isp1362_hc_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_017:sink_ready -> ISP1362_hc_translator_avalon_universal_slave_0_agent:rp_ready
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket                                    : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_018:sink_endofpacket
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rp_valid                                          : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_018:sink_valid
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket                                  : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_018:sink_startofpacket
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rp_data                                           : std_logic_vector(101 downto 0); -- ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_data -> id_router_018:sink_data
	signal isp1362_dc_translator_avalon_universal_slave_0_agent_rp_ready                                          : std_logic;                      -- id_router_018:sink_ready -> ISP1362_dc_translator_avalon_universal_slave_0_agent:rp_ready
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_019:sink_endofpacket
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_019:sink_valid
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_019:sink_startofpacket
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(101 downto 0); -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_019:sink_data
	signal audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_019:sink_ready -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                          : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_020:sink_endofpacket
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                                : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_020:sink_valid
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                        : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_020:sink_startofpacket
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                                 : std_logic_vector(101 downto 0); -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_020:sink_data
	signal vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                                : std_logic;                      -- id_router_020:sink_ready -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                        : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_021:sink_endofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                              : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_021:sink_valid
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                      : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_021:sink_startofpacket
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                               : std_logic_vector(101 downto 0); -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_021:sink_data
	signal dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                              : std_logic;                      -- id_router_021:sink_ready -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_022:sink_endofpacket
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_022:sink_valid
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_022:sink_startofpacket
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(101 downto 0); -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_022:sink_data
	signal seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                      -- id_router_022:sink_ready -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                         : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_023:sink_endofpacket
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                               : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_023:sink_valid
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                       : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_023:sink_startofpacket
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                                : std_logic_vector(83 downto 0);  -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_023:sink_data
	signal sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                               : std_logic;                      -- id_router_023:sink_ready -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket                   : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_024:sink_endofpacket
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                         : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_024:sink_valid
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket                 : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_024:sink_startofpacket
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                          : std_logic_vector(101 downto 0); -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_024:sink_data
	signal lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                         : std_logic;                      -- id_router_024:sink_ready -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                   : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_025:sink_endofpacket
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_valid                                         : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_025:sink_valid
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                 : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_025:sink_startofpacket
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_data                                          : std_logic_vector(101 downto 0); -- motor_cw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_025:sink_data
	signal motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_ready                                         : std_logic;                      -- id_router_025:sink_ready -> motor_cw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                  : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_026:sink_endofpacket
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_valid                                        : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_026:sink_valid
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                                : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_026:sink_startofpacket
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_data                                         : std_logic_vector(101 downto 0); -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_026:sink_data
	signal motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_ready                                        : std_logic;                      -- id_router_026:sink_ready -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal addr_router_src_endofpacket                                                                            : std_logic;                      -- addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	signal addr_router_src_valid                                                                                  : std_logic;                      -- addr_router:src_valid -> limiter:cmd_sink_valid
	signal addr_router_src_startofpacket                                                                          : std_logic;                      -- addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	signal addr_router_src_data                                                                                   : std_logic_vector(101 downto 0); -- addr_router:src_data -> limiter:cmd_sink_data
	signal addr_router_src_channel                                                                                : std_logic_vector(26 downto 0);  -- addr_router:src_channel -> limiter:cmd_sink_channel
	signal addr_router_src_ready                                                                                  : std_logic;                      -- limiter:cmd_sink_ready -> addr_router:src_ready
	signal limiter_rsp_src_endofpacket                                                                            : std_logic;                      -- limiter:rsp_src_endofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal limiter_rsp_src_valid                                                                                  : std_logic;                      -- limiter:rsp_src_valid -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal limiter_rsp_src_startofpacket                                                                          : std_logic;                      -- limiter:rsp_src_startofpacket -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal limiter_rsp_src_data                                                                                   : std_logic_vector(101 downto 0); -- limiter:rsp_src_data -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal limiter_rsp_src_channel                                                                                : std_logic_vector(26 downto 0);  -- limiter:rsp_src_channel -> cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal limiter_rsp_src_ready                                                                                  : std_logic;                      -- cpu_0_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	signal burst_adapter_source0_endofpacket                                                                      : std_logic;                      -- burst_adapter:source0_endofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_source0_valid                                                                            : std_logic;                      -- burst_adapter:source0_valid -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_source0_startofpacket                                                                    : std_logic;                      -- burst_adapter:source0_startofpacket -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_source0_data                                                                             : std_logic_vector(83 downto 0);  -- burst_adapter:source0_data -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_source0_ready                                                                            : std_logic;                      -- sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	signal burst_adapter_source0_channel                                                                          : std_logic_vector(26 downto 0);  -- burst_adapter:source0_channel -> sdram_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_001_source0_endofpacket                                                                  : std_logic;                      -- burst_adapter_001:source0_endofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_001_source0_valid                                                                        : std_logic;                      -- burst_adapter_001:source0_valid -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_001_source0_startofpacket                                                                : std_logic;                      -- burst_adapter_001:source0_startofpacket -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_001_source0_data                                                                         : std_logic_vector(74 downto 0);  -- burst_adapter_001:source0_data -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_001_source0_ready                                                                        : std_logic;                      -- cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	signal burst_adapter_001_source0_channel                                                                      : std_logic_vector(26 downto 0);  -- burst_adapter_001:source0_channel -> cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:cp_channel
	signal burst_adapter_002_source0_endofpacket                                                                  : std_logic;                      -- burst_adapter_002:source0_endofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal burst_adapter_002_source0_valid                                                                        : std_logic;                      -- burst_adapter_002:source0_valid -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal burst_adapter_002_source0_startofpacket                                                                : std_logic;                      -- burst_adapter_002:source0_startofpacket -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal burst_adapter_002_source0_data                                                                         : std_logic_vector(83 downto 0);  -- burst_adapter_002:source0_data -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal burst_adapter_002_source0_ready                                                                        : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	signal burst_adapter_002_source0_channel                                                                      : std_logic_vector(26 downto 0);  -- burst_adapter_002:source0_channel -> sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cpu_0_jtag_debug_module_reset_reset                                                                    : std_logic;                      -- cpu_0:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in0]
	signal rst_controller_001_reset_out_reset                                                                     : std_logic;                      -- rst_controller_001:reset_out -> [ISP1362_dc_translator:reset, ISP1362_dc_translator_avalon_universal_slave_0_agent:reset, ISP1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, ISP1362_hc_translator:reset, ISP1362_hc_translator_avalon_universal_slave_0_agent:reset, ISP1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_CLK_s1_translator:reset, SD_CLK_s1_translator_avalon_universal_slave_0_agent:reset, SD_CLK_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_CMD_s1_translator:reset, SD_CMD_s1_translator_avalon_universal_slave_0_agent:reset, SD_CMD_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SD_DAT_s1_translator:reset, SD_DAT_s1_translator_avalon_universal_slave_0_agent:reset, SD_DAT_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, addr_router:reset, addr_router_001:reset, burst_adapter:reset, burst_adapter_001:reset, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cfi_flash_0:reset_reset, cfi_flash_0_uas_translator:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cpu_0_data_master_translator:reset, cpu_0_data_master_translator_avalon_universal_master_0_agent:reset, cpu_0_instruction_master_translator:reset, cpu_0_instruction_master_translator_avalon_universal_master_0_agent:reset, cpu_0_jtag_debug_module_translator:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:reset, cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, epcs_controller_epcs_control_port_translator:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:reset, epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, id_router_007:reset, id_router_008:reset, id_router_009:reset, id_router_010:reset, id_router_011:reset, id_router_012:reset, id_router_013:reset, id_router_014:reset, id_router_015:reset, id_router_016:reset, id_router_017:reset, id_router_018:reset, irq_mapper:reset, jtag_uart_0_avalon_jtag_slave_translator:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, lcd_16207_0_control_slave_translator:reset, lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:reset, lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_green_s1_translator:reset, led_green_s1_translator_avalon_universal_slave_0_agent:reset, led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_red_s1_translator:reset, led_red_s1_translator_avalon_universal_slave_0_agent:reset, led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, rsp_xbar_demux_009:reset, rsp_xbar_demux_010:reset, rsp_xbar_demux_011:reset, rsp_xbar_demux_012:reset, rsp_xbar_demux_013:reset, rsp_xbar_demux_014:reset, rsp_xbar_demux_015:reset, rsp_xbar_demux_016:reset, rsp_xbar_demux_017:reset, rsp_xbar_demux_018:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_001_reset_out_reset:in, sdram_0_s1_translator:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, switch_pio_s1_translator:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent:reset, switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, sysid_qsys_0_control_slave_translator:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:reset, sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_0_s1_translator:reset, timer_0_s1_translator_avalon_universal_slave_0_agent:reset, timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, timer_1_s1_translator:reset, timer_1_s1_translator_avalon_universal_slave_0_agent:reset, timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, tri_state_bridge_0_bridge_0:reset, tri_state_bridge_0_pinSharer_0:reset_reset, uart_0_s1_translator:reset, uart_0_s1_translator_avalon_universal_slave_0_agent:reset, uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset]
	signal rst_controller_002_reset_out_reset                                                                     : std_logic;                      -- rst_controller_002:reset_out -> [Audio_0_avalon_slave_0_translator:reset, Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, DM9000A_avalon_slave_0_translator:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, SEG7_Display_avalon_slave_0_translator:reset, SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, VGA_0_avalon_slave_0_translator:reset, VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter_002:reset, id_router_019:reset, id_router_020:reset, id_router_021:reset, id_router_022:reset, id_router_023:reset, id_router_024:reset, id_router_025:reset, id_router_026:reset, lab7_FINAL_0_avalon_slave_0_translator:reset, lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, motor_ccw_s1_translator:reset, motor_ccw_s1_translator_avalon_universal_slave_0_agent:reset, motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, motor_cw_s1_translator:reset, motor_cw_s1_translator_avalon_universal_slave_0_agent:reset, motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux_019:reset, rsp_xbar_demux_020:reset, rsp_xbar_demux_021:reset, rsp_xbar_demux_022:reset, rsp_xbar_demux_023:reset, rsp_xbar_demux_024:reset, rsp_xbar_demux_025:reset, rsp_xbar_demux_026:reset, rst_controller_002_reset_out_reset:in, sram_0_avalon_slave_0_translator:reset, sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_004:reset, width_adapter_005:reset]
	signal cmd_xbar_demux_src0_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                            : std_logic_vector(26 downto 0);  -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                              : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                            : std_logic_vector(26 downto 0);  -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                              : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_src2_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src2_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	signal cmd_xbar_demux_src2_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src2_valid -> cmd_xbar_mux_002:sink0_valid
	signal cmd_xbar_demux_src2_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src2_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	signal cmd_xbar_demux_src2_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src2_data -> cmd_xbar_mux_002:sink0_data
	signal cmd_xbar_demux_src2_channel                                                                            : std_logic_vector(26 downto 0);  -- cmd_xbar_demux:src2_channel -> cmd_xbar_mux_002:sink0_channel
	signal cmd_xbar_demux_src2_ready                                                                              : std_logic;                      -- cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux:src2_ready
	signal cmd_xbar_demux_src3_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src3_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	signal cmd_xbar_demux_src3_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src3_valid -> cmd_xbar_mux_003:sink0_valid
	signal cmd_xbar_demux_src3_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src3_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	signal cmd_xbar_demux_src3_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src3_data -> cmd_xbar_mux_003:sink0_data
	signal cmd_xbar_demux_src3_channel                                                                            : std_logic_vector(26 downto 0);  -- cmd_xbar_demux:src3_channel -> cmd_xbar_mux_003:sink0_channel
	signal cmd_xbar_demux_src3_ready                                                                              : std_logic;                      -- cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux:src3_ready
	signal cmd_xbar_demux_src4_endofpacket                                                                        : std_logic;                      -- cmd_xbar_demux:src4_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	signal cmd_xbar_demux_src4_valid                                                                              : std_logic;                      -- cmd_xbar_demux:src4_valid -> cmd_xbar_mux_004:sink0_valid
	signal cmd_xbar_demux_src4_startofpacket                                                                      : std_logic;                      -- cmd_xbar_demux:src4_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	signal cmd_xbar_demux_src4_data                                                                               : std_logic_vector(101 downto 0); -- cmd_xbar_demux:src4_data -> cmd_xbar_mux_004:sink0_data
	signal cmd_xbar_demux_src4_channel                                                                            : std_logic_vector(26 downto 0);  -- cmd_xbar_demux:src4_channel -> cmd_xbar_mux_004:sink0_channel
	signal cmd_xbar_demux_src4_ready                                                                              : std_logic;                      -- cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux:src4_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                          : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                          : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal cmd_xbar_demux_001_src2_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	signal cmd_xbar_demux_001_src2_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_002:sink1_valid
	signal cmd_xbar_demux_001_src2_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	signal cmd_xbar_demux_001_src2_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_002:sink1_data
	signal cmd_xbar_demux_001_src2_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_002:sink1_channel
	signal cmd_xbar_demux_001_src2_ready                                                                          : std_logic;                      -- cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_001:src2_ready
	signal cmd_xbar_demux_001_src3_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	signal cmd_xbar_demux_001_src3_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_003:sink1_valid
	signal cmd_xbar_demux_001_src3_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	signal cmd_xbar_demux_001_src3_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_003:sink1_data
	signal cmd_xbar_demux_001_src3_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_003:sink1_channel
	signal cmd_xbar_demux_001_src3_ready                                                                          : std_logic;                      -- cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_001:src3_ready
	signal cmd_xbar_demux_001_src4_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	signal cmd_xbar_demux_001_src4_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_004:sink1_valid
	signal cmd_xbar_demux_001_src4_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	signal cmd_xbar_demux_001_src4_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_004:sink1_data
	signal cmd_xbar_demux_001_src4_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_004:sink1_channel
	signal cmd_xbar_demux_001_src4_ready                                                                          : std_logic;                      -- cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_001:src4_ready
	signal cmd_xbar_demux_001_src5_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src5_endofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src5_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src5_valid -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src5_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src5_startofpacket -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src5_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src5_data -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src5_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src5_channel -> jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src6_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src6_endofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src6_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src6_valid -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src6_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src6_startofpacket -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src6_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src6_data -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src6_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src6_channel -> uart_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src7_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src7_endofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src7_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src7_valid -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src7_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src7_startofpacket -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src7_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src7_data -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src7_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src7_channel -> timer_0_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src8_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src8_endofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src8_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src8_valid -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src8_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src8_startofpacket -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src8_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src8_data -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src8_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src8_channel -> timer_1_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src9_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux_001:src9_endofpacket -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src9_valid                                                                          : std_logic;                      -- cmd_xbar_demux_001:src9_valid -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src9_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux_001:src9_startofpacket -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src9_data                                                                           : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src9_data -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src9_channel                                                                        : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src9_channel -> lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src10_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src10_endofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src10_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src10_valid -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src10_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src10_startofpacket -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src10_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src10_data -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src10_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src10_channel -> led_red_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src11_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src11_endofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src11_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src11_valid -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src11_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src11_startofpacket -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src11_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src11_data -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src11_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src11_channel -> led_green_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src12_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src12_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src12_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src12_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src12_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src12_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src12_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src12_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src12_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src12_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src13_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src13_endofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src13_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src13_valid -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src13_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src13_startofpacket -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src13_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src13_data -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src13_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src13_channel -> switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src14_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src14_endofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src14_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src14_valid -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src14_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src14_startofpacket -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src14_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src14_data -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src14_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src14_channel -> SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src15_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src15_endofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src15_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src15_valid -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src15_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src15_startofpacket -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src15_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src15_data -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src15_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src15_channel -> SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src16_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src16_endofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src16_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src16_valid -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src16_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src16_startofpacket -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src16_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src16_data -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src16_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src16_channel -> SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src17_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src17_endofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src17_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src17_valid -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src17_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src17_startofpacket -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src17_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src17_data -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src17_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src17_channel -> ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src18_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src18_endofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src18_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src18_valid -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src18_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src18_startofpacket -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src18_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src18_data -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src18_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src18_channel -> ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src19_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src19_endofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src19_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src19_valid -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src19_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src19_startofpacket -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src19_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src19_data -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src19_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src19_channel -> Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src20_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src20_endofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src20_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src20_valid -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src20_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src20_startofpacket -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src20_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src20_data -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src20_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src20_channel -> VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src21_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src21_endofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src21_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src21_valid -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src21_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src21_startofpacket -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src21_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src21_data -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src21_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src21_channel -> DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src22_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src22_endofpacket -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src22_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src22_valid -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src22_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src22_startofpacket -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src22_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src22_data -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src22_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src22_channel -> SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src23_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src23_endofpacket -> width_adapter_004:in_endofpacket
	signal cmd_xbar_demux_001_src23_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src23_valid -> width_adapter_004:in_valid
	signal cmd_xbar_demux_001_src23_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src23_startofpacket -> width_adapter_004:in_startofpacket
	signal cmd_xbar_demux_001_src23_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src23_data -> width_adapter_004:in_data
	signal cmd_xbar_demux_001_src23_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src23_channel -> width_adapter_004:in_channel
	signal cmd_xbar_demux_001_src24_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src24_endofpacket -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src24_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src24_valid -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src24_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src24_startofpacket -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src24_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src24_data -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src24_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src24_channel -> lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src25_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src25_endofpacket -> motor_cw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src25_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src25_valid -> motor_cw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src25_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src25_startofpacket -> motor_cw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src25_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src25_data -> motor_cw_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src25_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src25_channel -> motor_cw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_demux_001_src26_endofpacket                                                                   : std_logic;                      -- cmd_xbar_demux_001:src26_endofpacket -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_demux_001_src26_valid                                                                         : std_logic;                      -- cmd_xbar_demux_001:src26_valid -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_demux_001_src26_startofpacket                                                                 : std_logic;                      -- cmd_xbar_demux_001:src26_startofpacket -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_demux_001_src26_data                                                                          : std_logic_vector(101 downto 0); -- cmd_xbar_demux_001:src26_data -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_demux_001_src26_channel                                                                       : std_logic_vector(26 downto 0);  -- cmd_xbar_demux_001:src26_channel -> motor_ccw_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal rsp_xbar_demux_src0_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                              : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                            : std_logic_vector(26 downto 0);  -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                              : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                        : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                              : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                      : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                               : std_logic_vector(101 downto 0); -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                            : std_logic_vector(26 downto 0);  -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                              : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_002_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	signal rsp_xbar_demux_002_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	signal rsp_xbar_demux_002_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	signal rsp_xbar_demux_002_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	signal rsp_xbar_demux_002_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	signal rsp_xbar_demux_002_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	signal rsp_xbar_demux_002_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	signal rsp_xbar_demux_002_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_001:sink2_valid
	signal rsp_xbar_demux_002_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	signal rsp_xbar_demux_002_src1_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_001:sink2_data
	signal rsp_xbar_demux_002_src1_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_001:sink2_channel
	signal rsp_xbar_demux_002_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_002:src1_ready
	signal rsp_xbar_demux_003_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	signal rsp_xbar_demux_003_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	signal rsp_xbar_demux_003_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	signal rsp_xbar_demux_003_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	signal rsp_xbar_demux_003_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	signal rsp_xbar_demux_003_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	signal rsp_xbar_demux_003_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	signal rsp_xbar_demux_003_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_001:sink3_valid
	signal rsp_xbar_demux_003_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	signal rsp_xbar_demux_003_src1_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_001:sink3_data
	signal rsp_xbar_demux_003_src1_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_001:sink3_channel
	signal rsp_xbar_demux_003_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_003:src1_ready
	signal rsp_xbar_demux_004_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux:sink4_endofpacket
	signal rsp_xbar_demux_004_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux:sink4_valid
	signal rsp_xbar_demux_004_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux:sink4_startofpacket
	signal rsp_xbar_demux_004_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_004:src0_data -> rsp_xbar_mux:sink4_data
	signal rsp_xbar_demux_004_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux:sink4_channel
	signal rsp_xbar_demux_004_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink4_ready -> rsp_xbar_demux_004:src0_ready
	signal rsp_xbar_demux_004_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	signal rsp_xbar_demux_004_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_001:sink4_valid
	signal rsp_xbar_demux_004_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	signal rsp_xbar_demux_004_src1_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_001:sink4_data
	signal rsp_xbar_demux_004_src1_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_001:sink4_channel
	signal rsp_xbar_demux_004_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_004:src1_ready
	signal rsp_xbar_demux_005_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	signal rsp_xbar_demux_005_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink5_valid
	signal rsp_xbar_demux_005_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	signal rsp_xbar_demux_005_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink5_data
	signal rsp_xbar_demux_005_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink5_channel
	signal rsp_xbar_demux_005_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink5_ready -> rsp_xbar_demux_005:src0_ready
	signal rsp_xbar_demux_006_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	signal rsp_xbar_demux_006_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink6_valid
	signal rsp_xbar_demux_006_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	signal rsp_xbar_demux_006_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink6_data
	signal rsp_xbar_demux_006_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink6_channel
	signal rsp_xbar_demux_006_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink6_ready -> rsp_xbar_demux_006:src0_ready
	signal rsp_xbar_demux_007_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_007:src0_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	signal rsp_xbar_demux_007_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_007:src0_valid -> rsp_xbar_mux_001:sink7_valid
	signal rsp_xbar_demux_007_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_007:src0_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	signal rsp_xbar_demux_007_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_007:src0_data -> rsp_xbar_mux_001:sink7_data
	signal rsp_xbar_demux_007_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_007:src0_channel -> rsp_xbar_mux_001:sink7_channel
	signal rsp_xbar_demux_007_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink7_ready -> rsp_xbar_demux_007:src0_ready
	signal rsp_xbar_demux_008_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_008:src0_endofpacket -> rsp_xbar_mux_001:sink8_endofpacket
	signal rsp_xbar_demux_008_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_008:src0_valid -> rsp_xbar_mux_001:sink8_valid
	signal rsp_xbar_demux_008_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_008:src0_startofpacket -> rsp_xbar_mux_001:sink8_startofpacket
	signal rsp_xbar_demux_008_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_008:src0_data -> rsp_xbar_mux_001:sink8_data
	signal rsp_xbar_demux_008_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_008:src0_channel -> rsp_xbar_mux_001:sink8_channel
	signal rsp_xbar_demux_008_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink8_ready -> rsp_xbar_demux_008:src0_ready
	signal rsp_xbar_demux_009_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_009:src0_endofpacket -> rsp_xbar_mux_001:sink9_endofpacket
	signal rsp_xbar_demux_009_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_009:src0_valid -> rsp_xbar_mux_001:sink9_valid
	signal rsp_xbar_demux_009_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_009:src0_startofpacket -> rsp_xbar_mux_001:sink9_startofpacket
	signal rsp_xbar_demux_009_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_009:src0_data -> rsp_xbar_mux_001:sink9_data
	signal rsp_xbar_demux_009_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_009:src0_channel -> rsp_xbar_mux_001:sink9_channel
	signal rsp_xbar_demux_009_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink9_ready -> rsp_xbar_demux_009:src0_ready
	signal rsp_xbar_demux_010_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_010:src0_endofpacket -> rsp_xbar_mux_001:sink10_endofpacket
	signal rsp_xbar_demux_010_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_010:src0_valid -> rsp_xbar_mux_001:sink10_valid
	signal rsp_xbar_demux_010_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_010:src0_startofpacket -> rsp_xbar_mux_001:sink10_startofpacket
	signal rsp_xbar_demux_010_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_010:src0_data -> rsp_xbar_mux_001:sink10_data
	signal rsp_xbar_demux_010_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_010:src0_channel -> rsp_xbar_mux_001:sink10_channel
	signal rsp_xbar_demux_010_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink10_ready -> rsp_xbar_demux_010:src0_ready
	signal rsp_xbar_demux_011_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_011:src0_endofpacket -> rsp_xbar_mux_001:sink11_endofpacket
	signal rsp_xbar_demux_011_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_011:src0_valid -> rsp_xbar_mux_001:sink11_valid
	signal rsp_xbar_demux_011_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_011:src0_startofpacket -> rsp_xbar_mux_001:sink11_startofpacket
	signal rsp_xbar_demux_011_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_011:src0_data -> rsp_xbar_mux_001:sink11_data
	signal rsp_xbar_demux_011_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_011:src0_channel -> rsp_xbar_mux_001:sink11_channel
	signal rsp_xbar_demux_011_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink11_ready -> rsp_xbar_demux_011:src0_ready
	signal rsp_xbar_demux_012_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_012:src0_endofpacket -> rsp_xbar_mux_001:sink12_endofpacket
	signal rsp_xbar_demux_012_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_012:src0_valid -> rsp_xbar_mux_001:sink12_valid
	signal rsp_xbar_demux_012_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_012:src0_startofpacket -> rsp_xbar_mux_001:sink12_startofpacket
	signal rsp_xbar_demux_012_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_012:src0_data -> rsp_xbar_mux_001:sink12_data
	signal rsp_xbar_demux_012_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_012:src0_channel -> rsp_xbar_mux_001:sink12_channel
	signal rsp_xbar_demux_012_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink12_ready -> rsp_xbar_demux_012:src0_ready
	signal rsp_xbar_demux_013_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_013:src0_endofpacket -> rsp_xbar_mux_001:sink13_endofpacket
	signal rsp_xbar_demux_013_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_013:src0_valid -> rsp_xbar_mux_001:sink13_valid
	signal rsp_xbar_demux_013_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_013:src0_startofpacket -> rsp_xbar_mux_001:sink13_startofpacket
	signal rsp_xbar_demux_013_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_013:src0_data -> rsp_xbar_mux_001:sink13_data
	signal rsp_xbar_demux_013_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_013:src0_channel -> rsp_xbar_mux_001:sink13_channel
	signal rsp_xbar_demux_013_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink13_ready -> rsp_xbar_demux_013:src0_ready
	signal rsp_xbar_demux_014_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_014:src0_endofpacket -> rsp_xbar_mux_001:sink14_endofpacket
	signal rsp_xbar_demux_014_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_014:src0_valid -> rsp_xbar_mux_001:sink14_valid
	signal rsp_xbar_demux_014_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_014:src0_startofpacket -> rsp_xbar_mux_001:sink14_startofpacket
	signal rsp_xbar_demux_014_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_014:src0_data -> rsp_xbar_mux_001:sink14_data
	signal rsp_xbar_demux_014_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_014:src0_channel -> rsp_xbar_mux_001:sink14_channel
	signal rsp_xbar_demux_014_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink14_ready -> rsp_xbar_demux_014:src0_ready
	signal rsp_xbar_demux_015_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_015:src0_endofpacket -> rsp_xbar_mux_001:sink15_endofpacket
	signal rsp_xbar_demux_015_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_015:src0_valid -> rsp_xbar_mux_001:sink15_valid
	signal rsp_xbar_demux_015_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_015:src0_startofpacket -> rsp_xbar_mux_001:sink15_startofpacket
	signal rsp_xbar_demux_015_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_015:src0_data -> rsp_xbar_mux_001:sink15_data
	signal rsp_xbar_demux_015_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_015:src0_channel -> rsp_xbar_mux_001:sink15_channel
	signal rsp_xbar_demux_015_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink15_ready -> rsp_xbar_demux_015:src0_ready
	signal rsp_xbar_demux_016_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_016:src0_endofpacket -> rsp_xbar_mux_001:sink16_endofpacket
	signal rsp_xbar_demux_016_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_016:src0_valid -> rsp_xbar_mux_001:sink16_valid
	signal rsp_xbar_demux_016_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_016:src0_startofpacket -> rsp_xbar_mux_001:sink16_startofpacket
	signal rsp_xbar_demux_016_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_016:src0_data -> rsp_xbar_mux_001:sink16_data
	signal rsp_xbar_demux_016_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_016:src0_channel -> rsp_xbar_mux_001:sink16_channel
	signal rsp_xbar_demux_016_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink16_ready -> rsp_xbar_demux_016:src0_ready
	signal rsp_xbar_demux_017_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_017:src0_endofpacket -> rsp_xbar_mux_001:sink17_endofpacket
	signal rsp_xbar_demux_017_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_017:src0_valid -> rsp_xbar_mux_001:sink17_valid
	signal rsp_xbar_demux_017_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_017:src0_startofpacket -> rsp_xbar_mux_001:sink17_startofpacket
	signal rsp_xbar_demux_017_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_017:src0_data -> rsp_xbar_mux_001:sink17_data
	signal rsp_xbar_demux_017_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_017:src0_channel -> rsp_xbar_mux_001:sink17_channel
	signal rsp_xbar_demux_017_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink17_ready -> rsp_xbar_demux_017:src0_ready
	signal rsp_xbar_demux_018_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_018:src0_endofpacket -> rsp_xbar_mux_001:sink18_endofpacket
	signal rsp_xbar_demux_018_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_018:src0_valid -> rsp_xbar_mux_001:sink18_valid
	signal rsp_xbar_demux_018_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_018:src0_startofpacket -> rsp_xbar_mux_001:sink18_startofpacket
	signal rsp_xbar_demux_018_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_018:src0_data -> rsp_xbar_mux_001:sink18_data
	signal rsp_xbar_demux_018_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_018:src0_channel -> rsp_xbar_mux_001:sink18_channel
	signal rsp_xbar_demux_018_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink18_ready -> rsp_xbar_demux_018:src0_ready
	signal rsp_xbar_demux_019_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_019:src0_endofpacket -> rsp_xbar_mux_001:sink19_endofpacket
	signal rsp_xbar_demux_019_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_019:src0_valid -> rsp_xbar_mux_001:sink19_valid
	signal rsp_xbar_demux_019_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_019:src0_startofpacket -> rsp_xbar_mux_001:sink19_startofpacket
	signal rsp_xbar_demux_019_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_019:src0_data -> rsp_xbar_mux_001:sink19_data
	signal rsp_xbar_demux_019_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_019:src0_channel -> rsp_xbar_mux_001:sink19_channel
	signal rsp_xbar_demux_019_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink19_ready -> rsp_xbar_demux_019:src0_ready
	signal rsp_xbar_demux_020_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_020:src0_endofpacket -> rsp_xbar_mux_001:sink20_endofpacket
	signal rsp_xbar_demux_020_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_020:src0_valid -> rsp_xbar_mux_001:sink20_valid
	signal rsp_xbar_demux_020_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_020:src0_startofpacket -> rsp_xbar_mux_001:sink20_startofpacket
	signal rsp_xbar_demux_020_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_020:src0_data -> rsp_xbar_mux_001:sink20_data
	signal rsp_xbar_demux_020_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_020:src0_channel -> rsp_xbar_mux_001:sink20_channel
	signal rsp_xbar_demux_020_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink20_ready -> rsp_xbar_demux_020:src0_ready
	signal rsp_xbar_demux_021_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_021:src0_endofpacket -> rsp_xbar_mux_001:sink21_endofpacket
	signal rsp_xbar_demux_021_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_021:src0_valid -> rsp_xbar_mux_001:sink21_valid
	signal rsp_xbar_demux_021_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_021:src0_startofpacket -> rsp_xbar_mux_001:sink21_startofpacket
	signal rsp_xbar_demux_021_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_021:src0_data -> rsp_xbar_mux_001:sink21_data
	signal rsp_xbar_demux_021_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_021:src0_channel -> rsp_xbar_mux_001:sink21_channel
	signal rsp_xbar_demux_021_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink21_ready -> rsp_xbar_demux_021:src0_ready
	signal rsp_xbar_demux_022_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_022:src0_endofpacket -> rsp_xbar_mux_001:sink22_endofpacket
	signal rsp_xbar_demux_022_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_022:src0_valid -> rsp_xbar_mux_001:sink22_valid
	signal rsp_xbar_demux_022_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_022:src0_startofpacket -> rsp_xbar_mux_001:sink22_startofpacket
	signal rsp_xbar_demux_022_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_022:src0_data -> rsp_xbar_mux_001:sink22_data
	signal rsp_xbar_demux_022_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_022:src0_channel -> rsp_xbar_mux_001:sink22_channel
	signal rsp_xbar_demux_022_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink22_ready -> rsp_xbar_demux_022:src0_ready
	signal rsp_xbar_demux_023_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_023:src0_endofpacket -> rsp_xbar_mux_001:sink23_endofpacket
	signal rsp_xbar_demux_023_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_023:src0_valid -> rsp_xbar_mux_001:sink23_valid
	signal rsp_xbar_demux_023_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_023:src0_startofpacket -> rsp_xbar_mux_001:sink23_startofpacket
	signal rsp_xbar_demux_023_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_023:src0_data -> rsp_xbar_mux_001:sink23_data
	signal rsp_xbar_demux_023_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_023:src0_channel -> rsp_xbar_mux_001:sink23_channel
	signal rsp_xbar_demux_023_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink23_ready -> rsp_xbar_demux_023:src0_ready
	signal rsp_xbar_demux_024_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_024:src0_endofpacket -> rsp_xbar_mux_001:sink24_endofpacket
	signal rsp_xbar_demux_024_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_024:src0_valid -> rsp_xbar_mux_001:sink24_valid
	signal rsp_xbar_demux_024_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_024:src0_startofpacket -> rsp_xbar_mux_001:sink24_startofpacket
	signal rsp_xbar_demux_024_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_024:src0_data -> rsp_xbar_mux_001:sink24_data
	signal rsp_xbar_demux_024_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_024:src0_channel -> rsp_xbar_mux_001:sink24_channel
	signal rsp_xbar_demux_024_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink24_ready -> rsp_xbar_demux_024:src0_ready
	signal rsp_xbar_demux_025_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_025:src0_endofpacket -> rsp_xbar_mux_001:sink25_endofpacket
	signal rsp_xbar_demux_025_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_025:src0_valid -> rsp_xbar_mux_001:sink25_valid
	signal rsp_xbar_demux_025_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_025:src0_startofpacket -> rsp_xbar_mux_001:sink25_startofpacket
	signal rsp_xbar_demux_025_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_025:src0_data -> rsp_xbar_mux_001:sink25_data
	signal rsp_xbar_demux_025_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_025:src0_channel -> rsp_xbar_mux_001:sink25_channel
	signal rsp_xbar_demux_025_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink25_ready -> rsp_xbar_demux_025:src0_ready
	signal rsp_xbar_demux_026_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux_026:src0_endofpacket -> rsp_xbar_mux_001:sink26_endofpacket
	signal rsp_xbar_demux_026_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux_026:src0_valid -> rsp_xbar_mux_001:sink26_valid
	signal rsp_xbar_demux_026_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux_026:src0_startofpacket -> rsp_xbar_mux_001:sink26_startofpacket
	signal rsp_xbar_demux_026_src0_data                                                                           : std_logic_vector(101 downto 0); -- rsp_xbar_demux_026:src0_data -> rsp_xbar_mux_001:sink26_data
	signal rsp_xbar_demux_026_src0_channel                                                                        : std_logic_vector(26 downto 0);  -- rsp_xbar_demux_026:src0_channel -> rsp_xbar_mux_001:sink26_channel
	signal rsp_xbar_demux_026_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink26_ready -> rsp_xbar_demux_026:src0_ready
	signal limiter_cmd_src_endofpacket                                                                            : std_logic;                      -- limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal limiter_cmd_src_startofpacket                                                                          : std_logic;                      -- limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal limiter_cmd_src_data                                                                                   : std_logic_vector(101 downto 0); -- limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	signal limiter_cmd_src_channel                                                                                : std_logic_vector(26 downto 0);  -- limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	signal limiter_cmd_src_ready                                                                                  : std_logic;                      -- cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                           : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	signal rsp_xbar_mux_src_valid                                                                                 : std_logic;                      -- rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	signal rsp_xbar_mux_src_startofpacket                                                                         : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	signal rsp_xbar_mux_src_data                                                                                  : std_logic_vector(101 downto 0); -- rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	signal rsp_xbar_mux_src_channel                                                                               : std_logic_vector(26 downto 0);  -- rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	signal rsp_xbar_mux_src_ready                                                                                 : std_logic;                      -- limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                        : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                              : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                      : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                               : std_logic_vector(101 downto 0); -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                            : std_logic_vector(26 downto 0);  -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                              : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                       : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                             : std_logic;                      -- rsp_xbar_mux_001:src_valid -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                     : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                              : std_logic_vector(101 downto 0); -- rsp_xbar_mux_001:src_data -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                           : std_logic_vector(26 downto 0);  -- rsp_xbar_mux_001:src_channel -> cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                             : std_logic;                      -- cpu_0_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                           : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_src_valid                                                                                 : std_logic;                      -- cmd_xbar_mux:src_valid -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_src_startofpacket                                                                         : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_src_data                                                                                  : std_logic_vector(101 downto 0); -- cmd_xbar_mux:src_data -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_src_channel                                                                               : std_logic_vector(26 downto 0);  -- cmd_xbar_mux:src_channel -> cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_src_ready                                                                                 : std_logic;                      -- cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux:src_ready
	signal id_router_src_endofpacket                                                                              : std_logic;                      -- id_router:src_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal id_router_src_valid                                                                                    : std_logic;                      -- id_router:src_valid -> rsp_xbar_demux:sink_valid
	signal id_router_src_startofpacket                                                                            : std_logic;                      -- id_router:src_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal id_router_src_data                                                                                     : std_logic_vector(101 downto 0); -- id_router:src_data -> rsp_xbar_demux:sink_data
	signal id_router_src_channel                                                                                  : std_logic_vector(26 downto 0);  -- id_router:src_channel -> rsp_xbar_demux:sink_channel
	signal id_router_src_ready                                                                                    : std_logic;                      -- rsp_xbar_demux:sink_ready -> id_router:src_ready
	signal cmd_xbar_mux_002_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_002:src_endofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_002_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_002:src_valid -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_002_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_002:src_startofpacket -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_002_src_data                                                                              : std_logic_vector(101 downto 0); -- cmd_xbar_mux_002:src_data -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_002_src_channel                                                                           : std_logic_vector(26 downto 0);  -- cmd_xbar_mux_002:src_channel -> epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_002_src_ready                                                                             : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_002:src_ready
	signal id_router_002_src_endofpacket                                                                          : std_logic;                      -- id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	signal id_router_002_src_valid                                                                                : std_logic;                      -- id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	signal id_router_002_src_startofpacket                                                                        : std_logic;                      -- id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	signal id_router_002_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	signal id_router_002_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	signal id_router_002_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	signal cmd_xbar_mux_004_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_004:src_endofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_004_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_004:src_valid -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_004_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_004:src_startofpacket -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_004_src_data                                                                              : std_logic_vector(101 downto 0); -- cmd_xbar_mux_004:src_data -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_004_src_channel                                                                           : std_logic_vector(26 downto 0);  -- cmd_xbar_mux_004:src_channel -> sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_004_src_ready                                                                             : std_logic;                      -- sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_004:src_ready
	signal id_router_004_src_endofpacket                                                                          : std_logic;                      -- id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	signal id_router_004_src_valid                                                                                : std_logic;                      -- id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	signal id_router_004_src_startofpacket                                                                        : std_logic;                      -- id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	signal id_router_004_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	signal id_router_004_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	signal id_router_004_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	signal cmd_xbar_demux_001_src5_ready                                                                          : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src5_ready
	signal id_router_005_src_endofpacket                                                                          : std_logic;                      -- id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	signal id_router_005_src_valid                                                                                : std_logic;                      -- id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	signal id_router_005_src_startofpacket                                                                        : std_logic;                      -- id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	signal id_router_005_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	signal id_router_005_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	signal id_router_005_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	signal cmd_xbar_demux_001_src6_ready                                                                          : std_logic;                      -- uart_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src6_ready
	signal id_router_006_src_endofpacket                                                                          : std_logic;                      -- id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	signal id_router_006_src_valid                                                                                : std_logic;                      -- id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	signal id_router_006_src_startofpacket                                                                        : std_logic;                      -- id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	signal id_router_006_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	signal id_router_006_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	signal id_router_006_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	signal cmd_xbar_demux_001_src7_ready                                                                          : std_logic;                      -- timer_0_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src7_ready
	signal id_router_007_src_endofpacket                                                                          : std_logic;                      -- id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	signal id_router_007_src_valid                                                                                : std_logic;                      -- id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	signal id_router_007_src_startofpacket                                                                        : std_logic;                      -- id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	signal id_router_007_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	signal id_router_007_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	signal id_router_007_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	signal cmd_xbar_demux_001_src8_ready                                                                          : std_logic;                      -- timer_1_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src8_ready
	signal id_router_008_src_endofpacket                                                                          : std_logic;                      -- id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	signal id_router_008_src_valid                                                                                : std_logic;                      -- id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	signal id_router_008_src_startofpacket                                                                        : std_logic;                      -- id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	signal id_router_008_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	signal id_router_008_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	signal id_router_008_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	signal cmd_xbar_demux_001_src9_ready                                                                          : std_logic;                      -- lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src9_ready
	signal id_router_009_src_endofpacket                                                                          : std_logic;                      -- id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	signal id_router_009_src_valid                                                                                : std_logic;                      -- id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	signal id_router_009_src_startofpacket                                                                        : std_logic;                      -- id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	signal id_router_009_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	signal id_router_009_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	signal id_router_009_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	signal cmd_xbar_demux_001_src10_ready                                                                         : std_logic;                      -- led_red_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src10_ready
	signal id_router_010_src_endofpacket                                                                          : std_logic;                      -- id_router_010:src_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	signal id_router_010_src_valid                                                                                : std_logic;                      -- id_router_010:src_valid -> rsp_xbar_demux_010:sink_valid
	signal id_router_010_src_startofpacket                                                                        : std_logic;                      -- id_router_010:src_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	signal id_router_010_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_010:src_data -> rsp_xbar_demux_010:sink_data
	signal id_router_010_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_010:src_channel -> rsp_xbar_demux_010:sink_channel
	signal id_router_010_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_010:sink_ready -> id_router_010:src_ready
	signal cmd_xbar_demux_001_src11_ready                                                                         : std_logic;                      -- led_green_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src11_ready
	signal id_router_011_src_endofpacket                                                                          : std_logic;                      -- id_router_011:src_endofpacket -> rsp_xbar_demux_011:sink_endofpacket
	signal id_router_011_src_valid                                                                                : std_logic;                      -- id_router_011:src_valid -> rsp_xbar_demux_011:sink_valid
	signal id_router_011_src_startofpacket                                                                        : std_logic;                      -- id_router_011:src_startofpacket -> rsp_xbar_demux_011:sink_startofpacket
	signal id_router_011_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_011:src_data -> rsp_xbar_demux_011:sink_data
	signal id_router_011_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_011:src_channel -> rsp_xbar_demux_011:sink_channel
	signal id_router_011_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_011:sink_ready -> id_router_011:src_ready
	signal cmd_xbar_demux_001_src12_ready                                                                         : std_logic;                      -- button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src12_ready
	signal id_router_012_src_endofpacket                                                                          : std_logic;                      -- id_router_012:src_endofpacket -> rsp_xbar_demux_012:sink_endofpacket
	signal id_router_012_src_valid                                                                                : std_logic;                      -- id_router_012:src_valid -> rsp_xbar_demux_012:sink_valid
	signal id_router_012_src_startofpacket                                                                        : std_logic;                      -- id_router_012:src_startofpacket -> rsp_xbar_demux_012:sink_startofpacket
	signal id_router_012_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_012:src_data -> rsp_xbar_demux_012:sink_data
	signal id_router_012_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_012:src_channel -> rsp_xbar_demux_012:sink_channel
	signal id_router_012_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_012:sink_ready -> id_router_012:src_ready
	signal cmd_xbar_demux_001_src13_ready                                                                         : std_logic;                      -- switch_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src13_ready
	signal id_router_013_src_endofpacket                                                                          : std_logic;                      -- id_router_013:src_endofpacket -> rsp_xbar_demux_013:sink_endofpacket
	signal id_router_013_src_valid                                                                                : std_logic;                      -- id_router_013:src_valid -> rsp_xbar_demux_013:sink_valid
	signal id_router_013_src_startofpacket                                                                        : std_logic;                      -- id_router_013:src_startofpacket -> rsp_xbar_demux_013:sink_startofpacket
	signal id_router_013_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_013:src_data -> rsp_xbar_demux_013:sink_data
	signal id_router_013_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_013:src_channel -> rsp_xbar_demux_013:sink_channel
	signal id_router_013_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_013:sink_ready -> id_router_013:src_ready
	signal cmd_xbar_demux_001_src14_ready                                                                         : std_logic;                      -- SD_DAT_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src14_ready
	signal id_router_014_src_endofpacket                                                                          : std_logic;                      -- id_router_014:src_endofpacket -> rsp_xbar_demux_014:sink_endofpacket
	signal id_router_014_src_valid                                                                                : std_logic;                      -- id_router_014:src_valid -> rsp_xbar_demux_014:sink_valid
	signal id_router_014_src_startofpacket                                                                        : std_logic;                      -- id_router_014:src_startofpacket -> rsp_xbar_demux_014:sink_startofpacket
	signal id_router_014_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_014:src_data -> rsp_xbar_demux_014:sink_data
	signal id_router_014_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_014:src_channel -> rsp_xbar_demux_014:sink_channel
	signal id_router_014_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_014:sink_ready -> id_router_014:src_ready
	signal cmd_xbar_demux_001_src15_ready                                                                         : std_logic;                      -- SD_CMD_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src15_ready
	signal id_router_015_src_endofpacket                                                                          : std_logic;                      -- id_router_015:src_endofpacket -> rsp_xbar_demux_015:sink_endofpacket
	signal id_router_015_src_valid                                                                                : std_logic;                      -- id_router_015:src_valid -> rsp_xbar_demux_015:sink_valid
	signal id_router_015_src_startofpacket                                                                        : std_logic;                      -- id_router_015:src_startofpacket -> rsp_xbar_demux_015:sink_startofpacket
	signal id_router_015_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_015:src_data -> rsp_xbar_demux_015:sink_data
	signal id_router_015_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_015:src_channel -> rsp_xbar_demux_015:sink_channel
	signal id_router_015_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_015:sink_ready -> id_router_015:src_ready
	signal cmd_xbar_demux_001_src16_ready                                                                         : std_logic;                      -- SD_CLK_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src16_ready
	signal id_router_016_src_endofpacket                                                                          : std_logic;                      -- id_router_016:src_endofpacket -> rsp_xbar_demux_016:sink_endofpacket
	signal id_router_016_src_valid                                                                                : std_logic;                      -- id_router_016:src_valid -> rsp_xbar_demux_016:sink_valid
	signal id_router_016_src_startofpacket                                                                        : std_logic;                      -- id_router_016:src_startofpacket -> rsp_xbar_demux_016:sink_startofpacket
	signal id_router_016_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_016:src_data -> rsp_xbar_demux_016:sink_data
	signal id_router_016_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_016:src_channel -> rsp_xbar_demux_016:sink_channel
	signal id_router_016_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_016:sink_ready -> id_router_016:src_ready
	signal cmd_xbar_demux_001_src17_ready                                                                         : std_logic;                      -- ISP1362_hc_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src17_ready
	signal id_router_017_src_endofpacket                                                                          : std_logic;                      -- id_router_017:src_endofpacket -> rsp_xbar_demux_017:sink_endofpacket
	signal id_router_017_src_valid                                                                                : std_logic;                      -- id_router_017:src_valid -> rsp_xbar_demux_017:sink_valid
	signal id_router_017_src_startofpacket                                                                        : std_logic;                      -- id_router_017:src_startofpacket -> rsp_xbar_demux_017:sink_startofpacket
	signal id_router_017_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_017:src_data -> rsp_xbar_demux_017:sink_data
	signal id_router_017_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_017:src_channel -> rsp_xbar_demux_017:sink_channel
	signal id_router_017_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_017:sink_ready -> id_router_017:src_ready
	signal cmd_xbar_demux_001_src18_ready                                                                         : std_logic;                      -- ISP1362_dc_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src18_ready
	signal id_router_018_src_endofpacket                                                                          : std_logic;                      -- id_router_018:src_endofpacket -> rsp_xbar_demux_018:sink_endofpacket
	signal id_router_018_src_valid                                                                                : std_logic;                      -- id_router_018:src_valid -> rsp_xbar_demux_018:sink_valid
	signal id_router_018_src_startofpacket                                                                        : std_logic;                      -- id_router_018:src_startofpacket -> rsp_xbar_demux_018:sink_startofpacket
	signal id_router_018_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_018:src_data -> rsp_xbar_demux_018:sink_data
	signal id_router_018_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_018:src_channel -> rsp_xbar_demux_018:sink_channel
	signal id_router_018_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_018:sink_ready -> id_router_018:src_ready
	signal cmd_xbar_demux_001_src19_ready                                                                         : std_logic;                      -- Audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src19_ready
	signal id_router_019_src_endofpacket                                                                          : std_logic;                      -- id_router_019:src_endofpacket -> rsp_xbar_demux_019:sink_endofpacket
	signal id_router_019_src_valid                                                                                : std_logic;                      -- id_router_019:src_valid -> rsp_xbar_demux_019:sink_valid
	signal id_router_019_src_startofpacket                                                                        : std_logic;                      -- id_router_019:src_startofpacket -> rsp_xbar_demux_019:sink_startofpacket
	signal id_router_019_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_019:src_data -> rsp_xbar_demux_019:sink_data
	signal id_router_019_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_019:src_channel -> rsp_xbar_demux_019:sink_channel
	signal id_router_019_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_019:sink_ready -> id_router_019:src_ready
	signal cmd_xbar_demux_001_src20_ready                                                                         : std_logic;                      -- VGA_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src20_ready
	signal id_router_020_src_endofpacket                                                                          : std_logic;                      -- id_router_020:src_endofpacket -> rsp_xbar_demux_020:sink_endofpacket
	signal id_router_020_src_valid                                                                                : std_logic;                      -- id_router_020:src_valid -> rsp_xbar_demux_020:sink_valid
	signal id_router_020_src_startofpacket                                                                        : std_logic;                      -- id_router_020:src_startofpacket -> rsp_xbar_demux_020:sink_startofpacket
	signal id_router_020_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_020:src_data -> rsp_xbar_demux_020:sink_data
	signal id_router_020_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_020:src_channel -> rsp_xbar_demux_020:sink_channel
	signal id_router_020_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_020:sink_ready -> id_router_020:src_ready
	signal cmd_xbar_demux_001_src21_ready                                                                         : std_logic;                      -- DM9000A_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src21_ready
	signal id_router_021_src_endofpacket                                                                          : std_logic;                      -- id_router_021:src_endofpacket -> rsp_xbar_demux_021:sink_endofpacket
	signal id_router_021_src_valid                                                                                : std_logic;                      -- id_router_021:src_valid -> rsp_xbar_demux_021:sink_valid
	signal id_router_021_src_startofpacket                                                                        : std_logic;                      -- id_router_021:src_startofpacket -> rsp_xbar_demux_021:sink_startofpacket
	signal id_router_021_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_021:src_data -> rsp_xbar_demux_021:sink_data
	signal id_router_021_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_021:src_channel -> rsp_xbar_demux_021:sink_channel
	signal id_router_021_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_021:sink_ready -> id_router_021:src_ready
	signal cmd_xbar_demux_001_src22_ready                                                                         : std_logic;                      -- SEG7_Display_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src22_ready
	signal id_router_022_src_endofpacket                                                                          : std_logic;                      -- id_router_022:src_endofpacket -> rsp_xbar_demux_022:sink_endofpacket
	signal id_router_022_src_valid                                                                                : std_logic;                      -- id_router_022:src_valid -> rsp_xbar_demux_022:sink_valid
	signal id_router_022_src_startofpacket                                                                        : std_logic;                      -- id_router_022:src_startofpacket -> rsp_xbar_demux_022:sink_startofpacket
	signal id_router_022_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_022:src_data -> rsp_xbar_demux_022:sink_data
	signal id_router_022_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_022:src_channel -> rsp_xbar_demux_022:sink_channel
	signal id_router_022_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_022:sink_ready -> id_router_022:src_ready
	signal cmd_xbar_demux_001_src24_ready                                                                         : std_logic;                      -- lab7_FINAL_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src24_ready
	signal id_router_024_src_endofpacket                                                                          : std_logic;                      -- id_router_024:src_endofpacket -> rsp_xbar_demux_024:sink_endofpacket
	signal id_router_024_src_valid                                                                                : std_logic;                      -- id_router_024:src_valid -> rsp_xbar_demux_024:sink_valid
	signal id_router_024_src_startofpacket                                                                        : std_logic;                      -- id_router_024:src_startofpacket -> rsp_xbar_demux_024:sink_startofpacket
	signal id_router_024_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_024:src_data -> rsp_xbar_demux_024:sink_data
	signal id_router_024_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_024:src_channel -> rsp_xbar_demux_024:sink_channel
	signal id_router_024_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_024:sink_ready -> id_router_024:src_ready
	signal cmd_xbar_demux_001_src25_ready                                                                         : std_logic;                      -- motor_cw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src25_ready
	signal id_router_025_src_endofpacket                                                                          : std_logic;                      -- id_router_025:src_endofpacket -> rsp_xbar_demux_025:sink_endofpacket
	signal id_router_025_src_valid                                                                                : std_logic;                      -- id_router_025:src_valid -> rsp_xbar_demux_025:sink_valid
	signal id_router_025_src_startofpacket                                                                        : std_logic;                      -- id_router_025:src_startofpacket -> rsp_xbar_demux_025:sink_startofpacket
	signal id_router_025_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_025:src_data -> rsp_xbar_demux_025:sink_data
	signal id_router_025_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_025:src_channel -> rsp_xbar_demux_025:sink_channel
	signal id_router_025_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_025:sink_ready -> id_router_025:src_ready
	signal cmd_xbar_demux_001_src26_ready                                                                         : std_logic;                      -- motor_ccw_s1_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux_001:src26_ready
	signal id_router_026_src_endofpacket                                                                          : std_logic;                      -- id_router_026:src_endofpacket -> rsp_xbar_demux_026:sink_endofpacket
	signal id_router_026_src_valid                                                                                : std_logic;                      -- id_router_026:src_valid -> rsp_xbar_demux_026:sink_valid
	signal id_router_026_src_startofpacket                                                                        : std_logic;                      -- id_router_026:src_startofpacket -> rsp_xbar_demux_026:sink_startofpacket
	signal id_router_026_src_data                                                                                 : std_logic_vector(101 downto 0); -- id_router_026:src_data -> rsp_xbar_demux_026:sink_data
	signal id_router_026_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_026:src_channel -> rsp_xbar_demux_026:sink_channel
	signal id_router_026_src_ready                                                                                : std_logic;                      -- rsp_xbar_demux_026:sink_ready -> id_router_026:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_001:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                              : std_logic_vector(101 downto 0); -- cmd_xbar_mux_001:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_001_src_channel                                                                           : std_logic_vector(26 downto 0);  -- cmd_xbar_mux_001:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_001_src_ready                                                                             : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux_001:src_ready
	signal width_adapter_src_endofpacket                                                                          : std_logic;                      -- width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	signal width_adapter_src_valid                                                                                : std_logic;                      -- width_adapter:out_valid -> burst_adapter:sink0_valid
	signal width_adapter_src_startofpacket                                                                        : std_logic;                      -- width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	signal width_adapter_src_data                                                                                 : std_logic_vector(83 downto 0);  -- width_adapter:out_data -> burst_adapter:sink0_data
	signal width_adapter_src_ready                                                                                : std_logic;                      -- burst_adapter:sink0_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                              : std_logic_vector(26 downto 0);  -- width_adapter:out_channel -> burst_adapter:sink0_channel
	signal id_router_001_src_endofpacket                                                                          : std_logic;                      -- id_router_001:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_001_src_valid                                                                                : std_logic;                      -- id_router_001:src_valid -> width_adapter_001:in_valid
	signal id_router_001_src_startofpacket                                                                        : std_logic;                      -- id_router_001:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_001_src_data                                                                                 : std_logic_vector(83 downto 0);  -- id_router_001:src_data -> width_adapter_001:in_data
	signal id_router_001_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_001:src_channel -> width_adapter_001:in_channel
	signal id_router_001_src_ready                                                                                : std_logic;                      -- width_adapter_001:in_ready -> id_router_001:src_ready
	signal width_adapter_001_src_endofpacket                                                                      : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal width_adapter_001_src_valid                                                                            : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux_001:sink_valid
	signal width_adapter_001_src_startofpacket                                                                    : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal width_adapter_001_src_data                                                                             : std_logic_vector(101 downto 0); -- width_adapter_001:out_data -> rsp_xbar_demux_001:sink_data
	signal width_adapter_001_src_ready                                                                            : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                          : std_logic_vector(26 downto 0);  -- width_adapter_001:out_channel -> rsp_xbar_demux_001:sink_channel
	signal cmd_xbar_mux_003_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux_003:src_endofpacket -> width_adapter_002:in_endofpacket
	signal cmd_xbar_mux_003_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux_003:src_valid -> width_adapter_002:in_valid
	signal cmd_xbar_mux_003_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux_003:src_startofpacket -> width_adapter_002:in_startofpacket
	signal cmd_xbar_mux_003_src_data                                                                              : std_logic_vector(101 downto 0); -- cmd_xbar_mux_003:src_data -> width_adapter_002:in_data
	signal cmd_xbar_mux_003_src_channel                                                                           : std_logic_vector(26 downto 0);  -- cmd_xbar_mux_003:src_channel -> width_adapter_002:in_channel
	signal cmd_xbar_mux_003_src_ready                                                                             : std_logic;                      -- width_adapter_002:in_ready -> cmd_xbar_mux_003:src_ready
	signal width_adapter_002_src_endofpacket                                                                      : std_logic;                      -- width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	signal width_adapter_002_src_valid                                                                            : std_logic;                      -- width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	signal width_adapter_002_src_startofpacket                                                                    : std_logic;                      -- width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	signal width_adapter_002_src_data                                                                             : std_logic_vector(74 downto 0);  -- width_adapter_002:out_data -> burst_adapter_001:sink0_data
	signal width_adapter_002_src_ready                                                                            : std_logic;                      -- burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	signal width_adapter_002_src_channel                                                                          : std_logic_vector(26 downto 0);  -- width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	signal id_router_003_src_endofpacket                                                                          : std_logic;                      -- id_router_003:src_endofpacket -> width_adapter_003:in_endofpacket
	signal id_router_003_src_valid                                                                                : std_logic;                      -- id_router_003:src_valid -> width_adapter_003:in_valid
	signal id_router_003_src_startofpacket                                                                        : std_logic;                      -- id_router_003:src_startofpacket -> width_adapter_003:in_startofpacket
	signal id_router_003_src_data                                                                                 : std_logic_vector(74 downto 0);  -- id_router_003:src_data -> width_adapter_003:in_data
	signal id_router_003_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_003:src_channel -> width_adapter_003:in_channel
	signal id_router_003_src_ready                                                                                : std_logic;                      -- width_adapter_003:in_ready -> id_router_003:src_ready
	signal width_adapter_003_src_endofpacket                                                                      : std_logic;                      -- width_adapter_003:out_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	signal width_adapter_003_src_valid                                                                            : std_logic;                      -- width_adapter_003:out_valid -> rsp_xbar_demux_003:sink_valid
	signal width_adapter_003_src_startofpacket                                                                    : std_logic;                      -- width_adapter_003:out_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	signal width_adapter_003_src_data                                                                             : std_logic_vector(101 downto 0); -- width_adapter_003:out_data -> rsp_xbar_demux_003:sink_data
	signal width_adapter_003_src_ready                                                                            : std_logic;                      -- rsp_xbar_demux_003:sink_ready -> width_adapter_003:out_ready
	signal width_adapter_003_src_channel                                                                          : std_logic_vector(26 downto 0);  -- width_adapter_003:out_channel -> rsp_xbar_demux_003:sink_channel
	signal cmd_xbar_demux_001_src23_ready                                                                         : std_logic;                      -- width_adapter_004:in_ready -> cmd_xbar_demux_001:src23_ready
	signal width_adapter_004_src_endofpacket                                                                      : std_logic;                      -- width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	signal width_adapter_004_src_valid                                                                            : std_logic;                      -- width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	signal width_adapter_004_src_startofpacket                                                                    : std_logic;                      -- width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	signal width_adapter_004_src_data                                                                             : std_logic_vector(83 downto 0);  -- width_adapter_004:out_data -> burst_adapter_002:sink0_data
	signal width_adapter_004_src_ready                                                                            : std_logic;                      -- burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	signal width_adapter_004_src_channel                                                                          : std_logic_vector(26 downto 0);  -- width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	signal id_router_023_src_endofpacket                                                                          : std_logic;                      -- id_router_023:src_endofpacket -> width_adapter_005:in_endofpacket
	signal id_router_023_src_valid                                                                                : std_logic;                      -- id_router_023:src_valid -> width_adapter_005:in_valid
	signal id_router_023_src_startofpacket                                                                        : std_logic;                      -- id_router_023:src_startofpacket -> width_adapter_005:in_startofpacket
	signal id_router_023_src_data                                                                                 : std_logic_vector(83 downto 0);  -- id_router_023:src_data -> width_adapter_005:in_data
	signal id_router_023_src_channel                                                                              : std_logic_vector(26 downto 0);  -- id_router_023:src_channel -> width_adapter_005:in_channel
	signal id_router_023_src_ready                                                                                : std_logic;                      -- width_adapter_005:in_ready -> id_router_023:src_ready
	signal width_adapter_005_src_endofpacket                                                                      : std_logic;                      -- width_adapter_005:out_endofpacket -> rsp_xbar_demux_023:sink_endofpacket
	signal width_adapter_005_src_valid                                                                            : std_logic;                      -- width_adapter_005:out_valid -> rsp_xbar_demux_023:sink_valid
	signal width_adapter_005_src_startofpacket                                                                    : std_logic;                      -- width_adapter_005:out_startofpacket -> rsp_xbar_demux_023:sink_startofpacket
	signal width_adapter_005_src_data                                                                             : std_logic_vector(101 downto 0); -- width_adapter_005:out_data -> rsp_xbar_demux_023:sink_data
	signal width_adapter_005_src_ready                                                                            : std_logic;                      -- rsp_xbar_demux_023:sink_ready -> width_adapter_005:out_ready
	signal width_adapter_005_src_channel                                                                          : std_logic_vector(26 downto 0);  -- width_adapter_005:out_channel -> rsp_xbar_demux_023:sink_channel
	signal limiter_cmd_valid_data                                                                                 : std_logic_vector(26 downto 0);  -- limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	signal irq_mapper_receiver0_irq                                                                               : std_logic;                      -- epcs_controller:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                                               : std_logic;                      -- jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                                               : std_logic;                      -- uart_0:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                                               : std_logic;                      -- timer_0:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                                               : std_logic;                      -- timer_1:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                                               : std_logic;                      -- button_pio:irq -> irq_mapper:receiver5_irq
	signal isp1362_hc_irq_irq                                                                                     : std_logic;                      -- ISP1362:avs_hc_irq_n_oINT0_N -> isp1362_hc_irq_irq:in
	signal isp1362_dc_irq_irq                                                                                     : std_logic;                      -- ISP1362:avs_dc_irq_n_oINT0_N -> isp1362_dc_irq_irq:in
	signal irq_mapper_receiver8_irq                                                                               : std_logic;                      -- DM9000A:oINT -> irq_mapper:receiver8_irq
	signal cpu_0_d_irq_irq                                                                                        : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> cpu_0:d_irq
	signal reset_n_ports_inv                                                                                      : std_logic;                      -- reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in1, rst_controller_002:reset_in0]
	signal sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- sdram_0_s1_translator_avalon_anti_slave_0_write:inv -> sdram_0:az_wr_n
	signal sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv                                               : std_logic;                      -- sdram_0_s1_translator_avalon_anti_slave_0_read:inv -> sdram_0:az_rd_n
	signal sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv                                         : std_logic_vector(1 downto 0);   -- sdram_0_s1_translator_avalon_anti_slave_0_byteenable:inv -> sdram_0:az_be_n
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write_ports_inv                       : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write:inv -> epcs_controller:write_n
	signal epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read_ports_inv                        : std_logic;                      -- epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read:inv -> epcs_controller:read_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv                           : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write:inv -> jtag_uart_0:av_write_n
	signal jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv                            : std_logic;                      -- jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read:inv -> jtag_uart_0:av_read_n
	signal uart_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                               : std_logic;                      -- uart_0_s1_translator_avalon_anti_slave_0_write:inv -> uart_0:write_n
	signal uart_0_s1_translator_avalon_anti_slave_0_read_ports_inv                                                : std_logic;                      -- uart_0_s1_translator_avalon_anti_slave_0_read:inv -> uart_0:read_n
	signal timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- timer_0_s1_translator_avalon_anti_slave_0_write:inv -> timer_0:write_n
	signal timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- timer_1_s1_translator_avalon_anti_slave_0_write:inv -> timer_1:write_n
	signal led_red_s1_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- led_red_s1_translator_avalon_anti_slave_0_write:inv -> led_red:write_n
	signal led_green_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                      -- led_green_s1_translator_avalon_anti_slave_0_write:inv -> led_green:write_n
	signal button_pio_s1_translator_avalon_anti_slave_0_write_ports_inv                                           : std_logic;                      -- button_pio_s1_translator_avalon_anti_slave_0_write:inv -> button_pio:write_n
	signal sd_dat_s1_translator_avalon_anti_slave_0_write_ports_inv                                               : std_logic;                      -- sd_dat_s1_translator_avalon_anti_slave_0_write:inv -> SD_DAT:write_n
	signal sd_cmd_s1_translator_avalon_anti_slave_0_write_ports_inv                                               : std_logic;                      -- sd_cmd_s1_translator_avalon_anti_slave_0_write:inv -> SD_CMD:write_n
	signal sd_clk_s1_translator_avalon_anti_slave_0_write_ports_inv                                               : std_logic;                      -- sd_clk_s1_translator_avalon_anti_slave_0_write:inv -> SD_CLK:write_n
	signal isp1362_hc_translator_avalon_anti_slave_0_chipselect_ports_inv                                         : std_logic;                      -- isp1362_hc_translator_avalon_anti_slave_0_chipselect:inv -> ISP1362:avs_hc_chipselect_n_iCS_N
	signal isp1362_hc_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- isp1362_hc_translator_avalon_anti_slave_0_write:inv -> ISP1362:avs_hc_write_n_iWR_N
	signal isp1362_hc_translator_avalon_anti_slave_0_read_ports_inv                                               : std_logic;                      -- isp1362_hc_translator_avalon_anti_slave_0_read:inv -> ISP1362:avs_hc_read_n_iRD_N
	signal isp1362_dc_translator_avalon_anti_slave_0_chipselect_ports_inv                                         : std_logic;                      -- isp1362_dc_translator_avalon_anti_slave_0_chipselect:inv -> ISP1362:avs_dc_chipselect_n_iCS_N
	signal isp1362_dc_translator_avalon_anti_slave_0_write_ports_inv                                              : std_logic;                      -- isp1362_dc_translator_avalon_anti_slave_0_write:inv -> ISP1362:avs_dc_write_n_iWR_N
	signal isp1362_dc_translator_avalon_anti_slave_0_read_ports_inv                                               : std_logic;                      -- isp1362_dc_translator_avalon_anti_slave_0_read:inv -> ISP1362:avs_dc_read_n_iRD_N
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv                             : std_logic;                      -- dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect:inv -> DM9000A:iCS_N
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv                                  : std_logic;                      -- dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write:inv -> DM9000A:iWR_N
	signal dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv                                   : std_logic;                      -- dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read:inv -> DM9000A:iRD_N
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv                              : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect:inv -> sram_0:iCE_N
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv                                   : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write:inv -> sram_0:iWE_N
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv                                    : std_logic;                      -- sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read:inv -> sram_0:iOE_N
	signal sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable_ports_inv                              : std_logic_vector(1 downto 0);   -- sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable:inv -> sram_0:iBE_N
	signal motor_cw_s1_translator_avalon_anti_slave_0_write_ports_inv                                             : std_logic;                      -- motor_cw_s1_translator_avalon_anti_slave_0_write:inv -> motor_cw:write_n
	signal motor_ccw_s1_translator_avalon_anti_slave_0_write_ports_inv                                            : std_logic;                      -- motor_ccw_s1_translator_avalon_anti_slave_0_write:inv -> motor_ccw:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                                                           : std_logic;                      -- rst_controller_001_reset_out_reset:inv -> [ISP1362:avs_dc_reset_n_iRST_N, ISP1362:avs_hc_reset_n_iRST_N, SD_CLK:reset_n, SD_CMD:reset_n, SD_DAT:reset_n, button_pio:reset_n, cpu_0:reset_n, epcs_controller:reset_n, jtag_uart_0:rst_n, lcd_16207_0:reset_n, led_green:reset_n, led_red:reset_n, sdram_0:reset_n, switch_pio:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, timer_1:reset_n, uart_0:reset_n]
	signal rst_controller_002_reset_out_reset_ports_inv                                                           : std_logic;                      -- rst_controller_002_reset_out_reset:inv -> [Audio_0:iRST_N, DM9000A:iRST_N, SEG7_Display:iRST_N, VGA_0:iRST_N, lab7_FINAL_0:resetn, motor_ccw:reset_n, motor_cw:reset_n, sram_0:iRST_N]
	signal irq_mapper_receiver6_inv                                                                               : std_logic;                      -- isp1362_hc_irq_irq:inv -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_inv                                                                               : std_logic;                      -- isp1362_dc_irq_irq:inv -> irq_mapper:receiver7_irq

begin

	sdram_0 : component system_0_sdram_0
		port map (
			clk            => clk_50,                                                         --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,                   -- reset.reset_n
			az_addr        => sdram_0_s1_translator_avalon_anti_slave_0_address,              --    s1.address
			az_be_n        => sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv, --      .byteenable_n
			az_cs          => sdram_0_s1_translator_avalon_anti_slave_0_chipselect,           --      .chipselect
			az_data        => sdram_0_s1_translator_avalon_anti_slave_0_writedata,            --      .writedata
			az_rd_n        => sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv,       --      .read_n
			az_wr_n        => sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv,      --      .write_n
			za_data        => sdram_0_s1_translator_avalon_anti_slave_0_readdata,             --      .readdata
			za_valid       => sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid,        --      .readdatavalid
			za_waitrequest => sdram_0_s1_translator_avalon_anti_slave_0_waitrequest,          --      .waitrequest
			zs_addr        => zs_addr_from_the_sdram_0,                                       --  wire.export
			zs_ba          => zs_ba_from_the_sdram_0,                                         --      .export
			zs_cas_n       => zs_cas_n_from_the_sdram_0,                                      --      .export
			zs_cke         => zs_cke_from_the_sdram_0,                                        --      .export
			zs_cs_n        => zs_cs_n_from_the_sdram_0,                                       --      .export
			zs_dq          => zs_dq_to_and_from_the_sdram_0,                                  --      .export
			zs_dqm         => zs_dqm_from_the_sdram_0,                                        --      .export
			zs_ras_n       => zs_ras_n_from_the_sdram_0,                                      --      .export
			zs_we_n        => zs_we_n_from_the_sdram_0                                        --      .export
		);

	epcs_controller : component system_0_epcs_controller
		port map (
			clk           => clk_50,                                                                           --               clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,                                     --             reset.reset_n
			address       => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address,         -- epcs_control_port.address
			chipselect    => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect,      --                  .chipselect
			dataavailable => open,                                                                             --                  .dataavailable
			endofpacket   => open,                                                                             --                  .endofpacket
			read_n        => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			readdata      => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			readyfordata  => open,                                                                             --                  .readyfordata
			write_n       => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			writedata     => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			irq           => irq_mapper_receiver0_irq                                                          --               irq.irq
		);

	jtag_uart_0 : component system_0_jtag_uart_0
		port map (
			clk            => clk_50,                                                                       --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                                 --             reset.reset_n
			av_chipselect  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address(0),      --                  .address
			av_read_n      => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv,  --                  .read_n
			av_readdata    => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,        --                  .readdata
			av_write_n     => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv, --                  .write_n
			av_writedata   => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,       --                  .writedata
			av_waitrequest => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                                      --               irq.irq
		);

	uart_0 : component system_0_uart_0
		port map (
			clk           => clk_50,                                                   --                 clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,             --               reset.reset_n
			address       => uart_0_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			begintransfer => uart_0_s1_translator_avalon_anti_slave_0_begintransfer,   --                    .begintransfer
			chipselect    => uart_0_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			read_n        => uart_0_s1_translator_avalon_anti_slave_0_read_ports_inv,  --                    .read_n
			write_n       => uart_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata     => uart_0_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			readdata      => uart_0_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			dataavailable => open,                                                     --                    .dataavailable
			readyfordata  => open,                                                     --                    .readyfordata
			rxd           => rxd_to_the_uart_0,                                        -- external_connection.export
			txd           => txd_from_the_uart_0,                                      --                    .export
			irq           => irq_mapper_receiver2_irq                                  --                 irq.irq
		);

	timer_0 : component system_0_timer_0
		port map (
			clk        => clk_50,                                                    --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,              -- reset.reset_n
			address    => timer_0_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_0_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_0_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_0_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver3_irq                                   --   irq.irq
		);

	timer_1 : component system_0_timer_0
		port map (
			clk        => clk_50,                                                    --   clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,              -- reset.reset_n
			address    => timer_1_s1_translator_avalon_anti_slave_0_address,         --    s1.address
			writedata  => timer_1_s1_translator_avalon_anti_slave_0_writedata,       --      .writedata
			readdata   => timer_1_s1_translator_avalon_anti_slave_0_readdata,        --      .readdata
			chipselect => timer_1_s1_translator_avalon_anti_slave_0_chipselect,      --      .chipselect
			write_n    => timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver4_irq                                   --   irq.irq
		);

	lcd_16207_0 : component system_0_lcd_16207_0
		port map (
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,                           --         reset.reset_n
			clk           => clk_50,                                                                 --           clk.clk
			begintransfer => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_begintransfer, -- control_slave.begintransfer
			read          => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_read,          --              .read
			write         => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_write,         --              .write
			readdata      => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_readdata,      --              .readdata
			writedata     => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_writedata,     --              .writedata
			address       => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_address,       --              .address
			LCD_RS        => LCD_RS_from_the_lcd_16207_0,                                            --      external.export
			LCD_RW        => LCD_RW_from_the_lcd_16207_0,                                            --              .export
			LCD_data      => LCD_data_to_and_from_the_lcd_16207_0,                                   --              .export
			LCD_E         => LCD_E_from_the_lcd_16207_0                                              --              .export
		);

	led_red : component system_0_led_red
		port map (
			clk        => clk_50,                                                    --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,              --               reset.reset_n
			address    => led_red_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_red_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_red_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_red_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_red_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => out_port_from_the_led_red                                  -- external_connection.export
		);

	led_green : component system_0_led_green
		port map (
			clk        => clk_50,                                                      --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => led_green_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => led_green_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => led_green_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => led_green_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => led_green_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => out_port_from_the_led_green                                  -- external_connection.export
		);

	button_pio : component system_0_button_pio
		port map (
			clk        => clk_50,                                                       --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,                 --               reset.reset_n
			address    => button_pio_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => button_pio_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => button_pio_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => button_pio_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => button_pio_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			in_port    => in_port_to_the_button_pio,                                    -- external_connection.export
			irq        => irq_mapper_receiver5_irq                                      --                 irq.irq
		);

	switch_pio : component system_0_switch_pio
		port map (
			clk      => clk_50,                                                --                 clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,          --               reset.reset_n
			address  => switch_pio_s1_translator_avalon_anti_slave_0_address,  --                  s1.address
			readdata => switch_pio_s1_translator_avalon_anti_slave_0_readdata, --                    .readdata
			in_port  => in_port_to_the_switch_pio                              -- external_connection.export
		);

	sd_dat : component system_0_SD_DAT
		port map (
			clk        => clk_50,                                                   --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => sd_dat_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => sd_dat_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => sd_dat_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => sd_dat_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => sd_dat_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			bidir_port => bidir_port_to_and_from_the_SD_DAT                         -- external_connection.export
		);

	sd_cmd : component system_0_SD_DAT
		port map (
			clk        => clk_50,                                                   --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => sd_cmd_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => sd_cmd_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => sd_cmd_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => sd_cmd_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => sd_cmd_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			bidir_port => bidir_port_to_and_from_the_SD_CMD                         -- external_connection.export
		);

	sd_clk : component system_0_SD_CLK
		port map (
			clk        => clk_50,                                                   --                 clk.clk
			reset_n    => rst_controller_001_reset_out_reset_ports_inv,             --               reset.reset_n
			address    => sd_clk_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => sd_clk_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => sd_clk_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => sd_clk_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => sd_clk_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => out_port_from_the_SD_CLK                                  -- external_connection.export
		);

	isp1362 : component ISP1362_IF
		port map (
			avs_hc_clk_iCLK           => clk_50,                                                         --    hc_clock.clk
			avs_hc_reset_n_iRST_N     => rst_controller_001_reset_out_reset_ports_inv,                   --  hc_reset_n.reset_n
			avs_hc_writedata_iDATA    => isp1362_hc_translator_avalon_anti_slave_0_writedata,            --          hc.writedata
			avs_hc_readdata_oDATA     => isp1362_hc_translator_avalon_anti_slave_0_readdata,             --            .readdata
			avs_hc_address_iADDR      => isp1362_hc_translator_avalon_anti_slave_0_address(0),           --            .address
			avs_hc_read_n_iRD_N       => isp1362_hc_translator_avalon_anti_slave_0_read_ports_inv,       --            .read_n
			avs_hc_write_n_iWR_N      => isp1362_hc_translator_avalon_anti_slave_0_write_ports_inv,      --            .write_n
			avs_hc_chipselect_n_iCS_N => isp1362_hc_translator_avalon_anti_slave_0_chipselect_ports_inv, --            .chipselect_n
			avs_hc_irq_n_oINT0_N      => isp1362_hc_irq_irq,                                             --      hc_irq.irq_n
			avs_dc_clk_iCLK           => clk_50,                                                         --    dc_clock.clk
			avs_dc_reset_n_iRST_N     => rst_controller_001_reset_out_reset_ports_inv,                   --  dc_reset_n.reset_n
			avs_dc_writedata_iDATA    => isp1362_dc_translator_avalon_anti_slave_0_writedata,            --          dc.writedata
			avs_dc_readdata_oDATA     => isp1362_dc_translator_avalon_anti_slave_0_readdata,             --            .readdata
			avs_dc_address_iADDR      => isp1362_dc_translator_avalon_anti_slave_0_address(0),           --            .address
			avs_dc_read_n_iRD_N       => isp1362_dc_translator_avalon_anti_slave_0_read_ports_inv,       --            .read_n
			avs_dc_write_n_iWR_N      => isp1362_dc_translator_avalon_anti_slave_0_write_ports_inv,      --            .write_n
			avs_dc_chipselect_n_iCS_N => isp1362_dc_translator_avalon_anti_slave_0_chipselect_ports_inv, --            .chipselect_n
			avs_dc_irq_n_oINT0_N      => isp1362_dc_irq_irq,                                             --      dc_irq.irq_n
			USB_DATA                  => USB_DATA_to_and_from_the_ISP1362,                               -- conduit_end.export
			USB_ADDR                  => USB_ADDR_from_the_ISP1362,                                      --            .export
			USB_RD_N                  => USB_RD_N_from_the_ISP1362,                                      --            .export
			USB_WR_N                  => USB_WR_N_from_the_ISP1362,                                      --            .export
			USB_CS_N                  => USB_CS_N_from_the_ISP1362,                                      --            .export
			USB_RST_N                 => USB_RST_N_from_the_ISP1362,                                     --            .export
			USB_INT0                  => USB_INT0_to_the_ISP1362,                                        --            .export
			USB_INT1                  => USB_INT1_to_the_ISP1362                                         --            .export
		);

	cpu_0 : component system_0_cpu_0
		port map (
			clk                                   => clk_50,                                                             --                       clk.clk
			reset_n                               => rst_controller_001_reset_out_reset_ports_inv,                       --                   reset_n.reset_n
			d_address                             => cpu_0_data_master_address,                                          --               data_master.address
			d_byteenable                          => cpu_0_data_master_byteenable,                                       --                          .byteenable
			d_read                                => cpu_0_data_master_read,                                             --                          .read
			d_readdata                            => cpu_0_data_master_readdata,                                         --                          .readdata
			d_waitrequest                         => cpu_0_data_master_waitrequest,                                      --                          .waitrequest
			d_write                               => cpu_0_data_master_write,                                            --                          .write
			d_writedata                           => cpu_0_data_master_writedata,                                        --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_0_data_master_debugaccess,                                      --                          .debugaccess
			i_address                             => cpu_0_instruction_master_address,                                   --        instruction_master.address
			i_read                                => cpu_0_instruction_master_read,                                      --                          .read
			i_readdata                            => cpu_0_instruction_master_readdata,                                  --                          .readdata
			i_waitrequest                         => cpu_0_instruction_master_waitrequest,                               --                          .waitrequest
			i_readdatavalid                       => cpu_0_instruction_master_readdatavalid,                             --                          .readdatavalid
			d_irq                                 => cpu_0_d_irq_irq,                                                    --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_0_jtag_debug_module_reset_reset,                                --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read,        --                          .read
			jtag_debug_module_readdata            => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write,       --                          .write
			jtag_debug_module_writedata           => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,   --                          .writedata
			no_ci_readra                          => open                                                                -- custom_instruction_master.readra
		);

	tri_state_bridge_0_bridge_0 : component system_0_tri_state_bridge_0_bridge_0
		port map (
			clk                               => clk_50,                                                             --   clk.clk
			reset                             => rst_controller_001_reset_out_reset,                                 -- reset.reset
			request                           => tri_state_bridge_0_pinsharer_0_tcm_request,                         --   tcs.request
			grant                             => tri_state_bridge_0_pinsharer_0_tcm_grant,                           --      .grant
			tcs_tri_state_bridge_0_data       => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out,     --      .tri_state_bridge_0_data_out
			tcs_tri_state_bridge_0_data_outen => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen,   --      .tri_state_bridge_0_data_outen
			tcs_tri_state_bridge_0_data_in    => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in,      --      .tri_state_bridge_0_data_in
			tcs_tri_state_bridge_0_readn      => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out,    --      .tri_state_bridge_0_readn_out
			tcs_write_n_to_the_cfi_flash_0    => tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out,  --      .write_n_to_the_cfi_flash_0_out
			tcs_tri_state_bridge_0_address    => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out,  --      .tri_state_bridge_0_address_out
			tcs_select_n_to_the_cfi_flash_0   => tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out, --      .select_n_to_the_cfi_flash_0_out
			tri_state_bridge_0_data           => tri_state_bridge_0_data,                                            --   out.tri_state_bridge_0_data
			tri_state_bridge_0_readn          => tri_state_bridge_0_readn,                                           --      .tri_state_bridge_0_readn
			write_n_to_the_cfi_flash_0        => write_n_to_the_cfi_flash_0,                                         --      .write_n_to_the_cfi_flash_0
			tri_state_bridge_0_address        => tri_state_bridge_0_address,                                         --      .tri_state_bridge_0_address
			select_n_to_the_cfi_flash_0       => select_n_to_the_cfi_flash_0                                         --      .select_n_to_the_cfi_flash_0
		);

	tri_state_bridge_0_pinsharer_0 : component system_0_tri_state_bridge_0_pinSharer_0
		port map (
			clk_clk                       => clk_50,                                                             --   clk.clk
			reset_reset                   => rst_controller_001_reset_out_reset,                                 -- reset.reset
			request                       => tri_state_bridge_0_pinsharer_0_tcm_request,                         --   tcm.request
			grant                         => tri_state_bridge_0_pinsharer_0_tcm_grant,                           --      .grant
			tri_state_bridge_0_address    => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_address_out,  --      .tri_state_bridge_0_address_out
			tri_state_bridge_0_readn      => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_readn_out,    --      .tri_state_bridge_0_readn_out
			write_n_to_the_cfi_flash_0    => tri_state_bridge_0_pinsharer_0_tcm_write_n_to_the_cfi_flash_0_out,  --      .write_n_to_the_cfi_flash_0_out
			tri_state_bridge_0_data       => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_out,     --      .tri_state_bridge_0_data_out
			tri_state_bridge_0_data_in    => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_in,      --      .tri_state_bridge_0_data_in
			tri_state_bridge_0_data_outen => tri_state_bridge_0_pinsharer_0_tcm_tri_state_bridge_0_data_outen,   --      .tri_state_bridge_0_data_outen
			select_n_to_the_cfi_flash_0   => tri_state_bridge_0_pinsharer_0_tcm_select_n_to_the_cfi_flash_0_out, --      .select_n_to_the_cfi_flash_0_out
			tcs0_request                  => cfi_flash_0_tcm_request,                                            --  tcs0.request
			tcs0_grant                    => cfi_flash_0_tcm_grant,                                              --      .grant
			tcs0_address_out              => cfi_flash_0_tcm_address_out,                                        --      .address_out
			tcs0_read_n_out(0)            => cfi_flash_0_tcm_read_n_out,                                         --      .read_n_out
			tcs0_write_n_out(0)           => cfi_flash_0_tcm_write_n_out,                                        --      .write_n_out
			tcs0_data_out                 => cfi_flash_0_tcm_data_out,                                           --      .data_out
			tcs0_data_in                  => cfi_flash_0_tcm_data_in,                                            --      .data_in
			tcs0_data_outen               => cfi_flash_0_tcm_data_outen,                                         --      .data_outen
			tcs0_chipselect_n_out(0)      => cfi_flash_0_tcm_chipselect_n_out                                    --      .chipselect_n_out
		);

	cfi_flash_0 : component system_0_cfi_flash_0
		generic map (
			TCM_ADDRESS_W                  => 22,
			TCM_DATA_W                     => 8,
			TCM_BYTEENABLE_W               => 1,
			TCM_READ_WAIT                  => 160,
			TCM_WRITE_WAIT                 => 160,
			TCM_SETUP_WAIT                 => 40,
			TCM_DATA_HOLD                  => 40,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 1,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 1,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 0,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 0,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 1,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 0,
			ACTIVE_LOW_OUTPUTENABLE        => 0,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk              => clk_50,                                                       --   clk.clk
			reset_reset          => rst_controller_001_reset_out_reset,                           -- reset.reset
			uas_address          => cfi_flash_0_uas_translator_avalon_anti_slave_0_address,       --   uas.address
			uas_burstcount       => cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount,    --      .burstcount
			uas_read             => cfi_flash_0_uas_translator_avalon_anti_slave_0_read,          --      .read
			uas_write            => cfi_flash_0_uas_translator_avalon_anti_slave_0_write,         --      .write
			uas_waitrequest      => cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest,   --      .waitrequest
			uas_readdatavalid    => cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid, --      .readdatavalid
			uas_byteenable       => cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable,    --      .byteenable
			uas_readdata         => cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata,      --      .readdata
			uas_writedata        => cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata,     --      .writedata
			uas_lock             => cfi_flash_0_uas_translator_avalon_anti_slave_0_lock,          --      .lock
			uas_debugaccess      => cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess,   --      .debugaccess
			tcm_write_n_out      => cfi_flash_0_tcm_write_n_out,                                  --   tcm.write_n_out
			tcm_read_n_out       => cfi_flash_0_tcm_read_n_out,                                   --      .read_n_out
			tcm_chipselect_n_out => cfi_flash_0_tcm_chipselect_n_out,                             --      .chipselect_n_out
			tcm_request          => cfi_flash_0_tcm_request,                                      --      .request
			tcm_grant            => cfi_flash_0_tcm_grant,                                        --      .grant
			tcm_address_out      => cfi_flash_0_tcm_address_out,                                  --      .address_out
			tcm_data_out         => cfi_flash_0_tcm_data_out,                                     --      .data_out
			tcm_data_outen       => cfi_flash_0_tcm_data_outen,                                   --      .data_outen
			tcm_data_in          => cfi_flash_0_tcm_data_in                                       --      .data_in
		);

	sysid_qsys_0 : component system_0_sysid_qsys_0
		port map (
			clock    => clk_50,                                                               --           clk.clk
			reset_n  => rst_controller_001_reset_out_reset_ports_inv,                         --         reset.reset_n
			readdata => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,   -- control_slave.readdata
			address  => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address(0)  --              .address
		);

	audio_0 : component AUDIO_DAC_FIFO
		generic map (
			REF_CLK     => 18432000,
			SAMPLE_RATE => 48000,
			DATA_WIDTH  => 16,
			CHANNEL_NUM => 2
		)
		port map (
			iWR_CLK   => clk_50,                                                          --                   clk.clk
			iRST_N    => rst_controller_002_reset_out_reset_ports_inv,                    --             clk_reset.reset_n
			oAUD_DATA => audio_0_oAUD_DATA,                                               -- avalon_slave_0_export.export
			oAUD_LRCK => audio_0_oAUD_LRCK,                                               --                      .export
			oAUD_BCK  => audio_0_oAUD_BCK,                                                --                      .export
			oAUD_XCK  => audio_0_oAUD_XCK,                                                --                      .export
			iCLK_18_4 => audio_0_iCLK_18_4,                                               --                      .export
			iDATA     => audio_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata, --        avalon_slave_0.writedata
			iWR       => audio_0_avalon_slave_0_translator_avalon_anti_slave_0_write,     --                      .write
			oDATA     => audio_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata   --                      .readdata
		);

	vga_0 : component VGA_NIOS_CTRL
		generic map (
			RAM_SIZE => 307200
		)
		port map (
			iCLK      => clk_50,                                                         --                   clk.clk
			iRST_N    => rst_controller_002_reset_out_reset_ports_inv,                   --             clk_reset.reset_n
			VGA_R     => vga_0_VGA_R,                                                    -- avalon_slave_0_export.export
			VGA_G     => vga_0_VGA_G,                                                    --                      .export
			VGA_B     => vga_0_VGA_B,                                                    --                      .export
			VGA_HS    => vga_0_VGA_HS,                                                   --                      .export
			VGA_VS    => vga_0_VGA_VS,                                                   --                      .export
			VGA_SYNC  => vga_0_VGA_SYNC,                                                 --                      .export
			VGA_BLANK => vga_0_VGA_BLANK,                                                --                      .export
			VGA_CLK   => vga_0_VGA_CLK,                                                  --                      .export
			iCLK_25   => vga_0_iCLK_25,                                                  --                      .export
			oDATA     => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,   --        avalon_slave_0.readdata
			iDATA     => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,  --                      .writedata
			iADDR     => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_address,    --                      .address
			iWR       => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_write,      --                      .write
			iRD       => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_read,       --                      .read
			iCS       => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect  --                      .chipselect
		);

	dm9000a : component DM9000A_IF
		port map (
			iCLK       => clk_50,                                                                     --                   clk.clk
			iRST_N     => rst_controller_002_reset_out_reset_ports_inv,                               --             clk_reset.reset_n
			iOSC_50    => dm9000a_iOSC_50,                                                            -- avalon_slave_0_export.export
			ENET_DATA  => dm9000a_ENET_DATA,                                                          --                      .export
			ENET_CMD   => dm9000a_ENET_CMD,                                                           --                      .export
			ENET_RD_N  => dm9000a_ENET_RD_N,                                                          --                      .export
			ENET_WR_N  => dm9000a_ENET_WR_N,                                                          --                      .export
			ENET_CS_N  => dm9000a_ENET_CS_N,                                                          --                      .export
			ENET_RST_N => dm9000a_ENET_RST_N,                                                         --                      .export
			ENET_CLK   => dm9000a_ENET_CLK,                                                           --                      .export
			ENET_INT   => dm9000a_ENET_INT,                                                           --                      .export
			iDATA      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata,            --        avalon_slave_0.writedata
			iCMD       => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address(0),           --                      .address
			iRD_N      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv,       --                      .read_n
			iWR_N      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv,      --                      .write_n
			iCS_N      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv, --                      .chipselect_n
			oDATA      => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata,             --                      .readdata
			oINT       => irq_mapper_receiver8_irq                                                    --    avalon_slave_0_irq.irq
		);

	seg7_display : component SEG7_LUT_8
		port map (
			iCLK   => clk_50,                                                               --                   clk.clk
			iRST_N => rst_controller_002_reset_out_reset_ports_inv,                         --             clk_reset.reset_n
			oSEG0  => seg7_display_oSEG0,                                                   -- avalon_slave_0_export.export
			oSEG1  => seg7_display_oSEG1,                                                   --                      .export
			oSEG2  => seg7_display_oSEG2,                                                   --                      .export
			oSEG3  => seg7_display_oSEG3,                                                   --                      .export
			oSEG4  => seg7_display_oSEG4,                                                   --                      .export
			oSEG5  => seg7_display_oSEG5,                                                   --                      .export
			oSEG6  => seg7_display_oSEG6,                                                   --                      .export
			oSEG7  => seg7_display_oSEG7,                                                   --                      .export
			iDIG   => seg7_display_avalon_slave_0_translator_avalon_anti_slave_0_writedata, --        avalon_slave_0.writedata
			iWR    => seg7_display_avalon_slave_0_translator_avalon_anti_slave_0_write      --                      .write
		);

	sram_0 : component SRAM_16Bit_512K
		port map (
			iCLK      => clk_50,                                                                    --                   clk.clk
			iRST_N    => rst_controller_002_reset_out_reset_ports_inv,                              --             clk_reset.reset_n
			SRAM_DQ   => sram_0_avalon_slave_0_export_DQ,                                           -- avalon_slave_0_export.export
			SRAM_ADDR => sram_0_avalon_slave_0_export_ADDR,                                         --                      .export
			SRAM_UB_N => sram_0_avalon_slave_0_export_UB_N,                                         --                      .export
			SRAM_LB_N => sram_0_avalon_slave_0_export_LB_N,                                         --                      .export
			SRAM_WE_N => sram_0_avalon_slave_0_export_WE_N,                                         --                      .export
			SRAM_CE_N => sram_0_avalon_slave_0_export_CE_N,                                         --                      .export
			SRAM_OE_N => sram_0_avalon_slave_0_export_OE_N,                                         --                      .export
			iDATA     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,            --        avalon_slave_0.writedata
			oDATA     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,             --                      .readdata
			iADDR     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address,              --                      .address
			iWE_N     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv,      --                      .write_n
			iOE_N     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv,       --                      .read_n
			iCE_N     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv, --                      .chipselect_n
			iBE_N     => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable_ports_inv  --                      .byteenable_n
		);

	lab7_final_0 : component top_avalon
		port map (
			chipselect => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect, -- avalon_slave_0.chipselect
			writedata  => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,  --               .writedata
			readdata   => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,   --               .readdata
			add        => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_address(0), --               .address
			write_en   => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write,      --               .write
			read_en    => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_read,       --               .read
			clock      => clk_50,                                                                --     clock_sink.clk
			resetn     => rst_controller_002_reset_out_reset_ports_inv                           --     reset_sink.reset_n
		);

	motor_cw : component system_0_SD_CLK
		port map (
			clk        => clk_50,                                                     --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,               --               reset.reset_n
			address    => motor_cw_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => motor_cw_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => motor_cw_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => motor_cw_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => motor_cw_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => cw_output_export                                            -- external_connection.export
		);

	motor_ccw : component system_0_SD_CLK
		port map (
			clk        => clk_50,                                                      --                 clk.clk
			reset_n    => rst_controller_002_reset_out_reset_ports_inv,                --               reset.reset_n
			address    => motor_ccw_s1_translator_avalon_anti_slave_0_address,         --                  s1.address
			write_n    => motor_ccw_s1_translator_avalon_anti_slave_0_write_ports_inv, --                    .write_n
			writedata  => motor_ccw_s1_translator_avalon_anti_slave_0_writedata,       --                    .writedata
			chipselect => motor_ccw_s1_translator_avalon_anti_slave_0_chipselect,      --                    .chipselect
			readdata   => motor_ccw_s1_translator_avalon_anti_slave_0_readdata,        --                    .readdata
			out_port   => ccw_output_export                                            -- external_connection.export
		);

	cpu_0_instruction_master_translator : component system_0_cpu_0_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 1,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_50,                                                                      --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                          --                     reset.reset
			uav_address              => cpu_0_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_0_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_0_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_0_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_0_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_0_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_0_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_0_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_0_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_0_instruction_master_readdata,                                           --                          .readdata
			av_readdatavalid         => cpu_0_instruction_master_readdatavalid,                                      --                          .readdatavalid
			av_burstcount            => "1",                                                                         --               (terminated)
			av_byteenable            => "1111",                                                                      --               (terminated)
			av_beginbursttransfer    => '0',                                                                         --               (terminated)
			av_begintransfer         => '0',                                                                         --               (terminated)
			av_chipselect            => '0',                                                                         --               (terminated)
			av_write                 => '0',                                                                         --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                          --               (terminated)
			av_lock                  => '0',                                                                         --               (terminated)
			av_debugaccess           => '0',                                                                         --               (terminated)
			uav_clken                => open,                                                                        --               (terminated)
			av_clken                 => '1',                                                                         --               (terminated)
			uav_response             => "00",                                                                        --               (terminated)
			av_response              => open,                                                                        --               (terminated)
			uav_writeresponserequest => open,                                                                        --               (terminated)
			uav_writeresponsevalid   => '0',                                                                         --               (terminated)
			av_writeresponserequest  => '0',                                                                         --               (terminated)
			av_writeresponsevalid    => open                                                                         --               (terminated)
		);

	cpu_0_data_master_translator : component system_0_cpu_0_data_master_translator
		generic map (
			AV_ADDRESS_W                => 25,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 25,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_50,                                                               --                       clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                   --                     reset.reset
			uav_address              => cpu_0_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_0_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_0_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_0_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_0_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_0_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_0_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_0_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_0_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_0_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_0_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_0_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_0_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_0_data_master_read,                                               --                          .read
			av_readdata              => cpu_0_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_0_data_master_write,                                              --                          .write
			av_writedata             => cpu_0_data_master_writedata,                                          --                          .writedata
			av_debugaccess           => cpu_0_data_master_debugaccess,                                        --                          .debugaccess
			av_burstcount            => "1",                                                                  --               (terminated)
			av_beginbursttransfer    => '0',                                                                  --               (terminated)
			av_begintransfer         => '0',                                                                  --               (terminated)
			av_chipselect            => '0',                                                                  --               (terminated)
			av_readdatavalid         => open,                                                                 --               (terminated)
			av_lock                  => '0',                                                                  --               (terminated)
			uav_clken                => open,                                                                 --               (terminated)
			av_clken                 => '1',                                                                  --               (terminated)
			uav_response             => "00",                                                                 --               (terminated)
			av_response              => open,                                                                 --               (terminated)
			uav_writeresponserequest => open,                                                                 --               (terminated)
			uav_writeresponsevalid   => '0',                                                                  --               (terminated)
			av_writeresponserequest  => '0',                                                                  --               (terminated)
			av_writeresponsevalid    => open                                                                  --               (terminated)
		);

	cpu_0_jtag_debug_module_translator : component system_0_cpu_0_jtag_debug_module_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                             --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                 --                    reset.reset
			uav_address              => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_waitrequest           => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_debugaccess           => cpu_0_jtag_debug_module_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                               --              (terminated)
			av_beginbursttransfer    => open,                                                                               --              (terminated)
			av_burstcount            => open,                                                                               --              (terminated)
			av_readdatavalid         => '0',                                                                                --              (terminated)
			av_writebyteenable       => open,                                                                               --              (terminated)
			av_lock                  => open,                                                                               --              (terminated)
			av_chipselect            => open,                                                                               --              (terminated)
			av_clken                 => open,                                                                               --              (terminated)
			uav_clken                => '0',                                                                                --              (terminated)
			av_outputenable          => open,                                                                               --              (terminated)
			uav_response             => open,                                                                               --              (terminated)
			av_response              => "00",                                                                               --              (terminated)
			uav_writeresponserequest => '0',                                                                                --              (terminated)
			uav_writeresponsevalid   => open,                                                                               --              (terminated)
			av_writeresponserequest  => open,                                                                               --              (terminated)
			av_writeresponsevalid    => '0'                                                                                 --              (terminated)
		);

	sdram_0_s1_translator : component system_0_sdram_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                    reset.reset
			uav_address              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sdram_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sdram_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sdram_0_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sdram_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sdram_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sdram_0_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => sdram_0_s1_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => sdram_0_s1_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => sdram_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	epcs_controller_epcs_control_port_translator : component system_0_epcs_controller_epcs_control_port_translator
		generic map (
			AV_ADDRESS_W                   => 9,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                                       --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                           --                    reset.reset
			uav_address              => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                         --              (terminated)
			av_beginbursttransfer    => open,                                                                                         --              (terminated)
			av_burstcount            => open,                                                                                         --              (terminated)
			av_byteenable            => open,                                                                                         --              (terminated)
			av_readdatavalid         => '0',                                                                                          --              (terminated)
			av_waitrequest           => '0',                                                                                          --              (terminated)
			av_writebyteenable       => open,                                                                                         --              (terminated)
			av_lock                  => open,                                                                                         --              (terminated)
			av_clken                 => open,                                                                                         --              (terminated)
			uav_clken                => '0',                                                                                          --              (terminated)
			av_debugaccess           => open,                                                                                         --              (terminated)
			av_outputenable          => open,                                                                                         --              (terminated)
			uav_response             => open,                                                                                         --              (terminated)
			av_response              => "00",                                                                                         --              (terminated)
			uav_writeresponserequest => '0',                                                                                          --              (terminated)
			uav_writeresponsevalid   => open,                                                                                         --              (terminated)
			av_writeresponserequest  => open,                                                                                         --              (terminated)
			av_writeresponsevalid    => '0'                                                                                           --              (terminated)
		);

	cfi_flash_0_uas_translator : component system_0_cfi_flash_0_uas_translator
		generic map (
			AV_ADDRESS_W                   => 22,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 8,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 1,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 1,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 1,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 1,
			AV_ADDRESS_SYMBOLS             => 1,
			AV_BURSTCOUNT_SYMBOLS          => 1,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                     --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                         --                    reset.reset
			uav_address              => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => cfi_flash_0_uas_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => cfi_flash_0_uas_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => cfi_flash_0_uas_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => cfi_flash_0_uas_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => cfi_flash_0_uas_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_burstcount            => cfi_flash_0_uas_translator_avalon_anti_slave_0_burstcount,                  --                         .burstcount
			av_byteenable            => cfi_flash_0_uas_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_readdatavalid         => cfi_flash_0_uas_translator_avalon_anti_slave_0_readdatavalid,               --                         .readdatavalid
			av_waitrequest           => cfi_flash_0_uas_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_lock                  => cfi_flash_0_uas_translator_avalon_anti_slave_0_lock,                        --                         .lock
			av_debugaccess           => cfi_flash_0_uas_translator_avalon_anti_slave_0_debugaccess,                 --                         .debugaccess
			av_begintransfer         => open,                                                                       --              (terminated)
			av_beginbursttransfer    => open,                                                                       --              (terminated)
			av_writebyteenable       => open,                                                                       --              (terminated)
			av_chipselect            => open,                                                                       --              (terminated)
			av_clken                 => open,                                                                       --              (terminated)
			uav_clken                => '0',                                                                        --              (terminated)
			av_outputenable          => open,                                                                       --              (terminated)
			uav_response             => open,                                                                       --              (terminated)
			av_response              => "00",                                                                       --              (terminated)
			uav_writeresponserequest => '0',                                                                        --              (terminated)
			uav_writeresponsevalid   => open,                                                                       --              (terminated)
			av_writeresponserequest  => open,                                                                       --              (terminated)
			av_writeresponsevalid    => '0'                                                                         --              (terminated)
		);

	sysid_qsys_0_control_slave_translator : component system_0_sysid_qsys_0_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                    --                    reset.reset
			uav_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => sysid_qsys_0_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                                  --              (terminated)
			av_read                  => open,                                                                                  --              (terminated)
			av_writedata             => open,                                                                                  --              (terminated)
			av_begintransfer         => open,                                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                                  --              (terminated)
			av_burstcount            => open,                                                                                  --              (terminated)
			av_byteenable            => open,                                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                                  --              (terminated)
			av_lock                  => open,                                                                                  --              (terminated)
			av_chipselect            => open,                                                                                  --              (terminated)
			av_clken                 => open,                                                                                  --              (terminated)
			uav_clken                => '0',                                                                                   --              (terminated)
			av_debugaccess           => open,                                                                                  --              (terminated)
			av_outputenable          => open,                                                                                  --              (terminated)
			uav_response             => open,                                                                                  --              (terminated)
			av_response              => "00",                                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                                    --              (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator : component system_0_jtag_uart_0_avalon_jtag_slave_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 1,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                                   --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                       --                    reset.reset
			uav_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_waitrequest           => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest,                 --                         .waitrequest
			av_chipselect            => jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                     --              (terminated)
			av_byteenable            => open,                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                     --              (terminated)
			av_lock                  => open,                                                                                     --              (terminated)
			av_clken                 => open,                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                     --              (terminated)
			uav_response             => open,                                                                                     --              (terminated)
			av_response              => "00",                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                       --              (terminated)
		);

	uart_0_s1_translator : component system_0_uart_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                   --                    reset.reset
			uav_address              => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => uart_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => uart_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => uart_0_s1_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => uart_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => uart_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => uart_0_s1_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_chipselect            => uart_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	timer_0_s1_translator : component system_0_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                    reset.reset
			uav_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_0_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_0_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_0_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_0_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_0_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	timer_1_s1_translator : component system_0_timer_0_s1_translator
		generic map (
			AV_ADDRESS_W                   => 3,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                    reset.reset
			uav_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => timer_1_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => timer_1_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => timer_1_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => timer_1_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => timer_1_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	lcd_16207_0_control_slave_translator : component system_0_lcd_16207_0_control_slave_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 8,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 13,
			AV_WRITE_WAIT_CYCLES           => 13,
			AV_SETUP_WAIT_CYCLES           => 13,
			AV_DATA_HOLD_CYCLES            => 13
		)
		port map (
			clk                      => clk_50,                                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                                   --                    reset.reset
			uav_address              => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_begintransfer         => lcd_16207_0_control_slave_translator_avalon_anti_slave_0_begintransfer,               --                         .begintransfer
			av_beginbursttransfer    => open,                                                                                 --              (terminated)
			av_burstcount            => open,                                                                                 --              (terminated)
			av_byteenable            => open,                                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                                 --              (terminated)
			av_lock                  => open,                                                                                 --              (terminated)
			av_chipselect            => open,                                                                                 --              (terminated)
			av_clken                 => open,                                                                                 --              (terminated)
			uav_clken                => '0',                                                                                  --              (terminated)
			av_debugaccess           => open,                                                                                 --              (terminated)
			av_outputenable          => open,                                                                                 --              (terminated)
			uav_response             => open,                                                                                 --              (terminated)
			av_response              => "00",                                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                                   --              (terminated)
		);

	led_red_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                    reset.reset
			uav_address              => led_red_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => led_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => led_red_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => led_red_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => led_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => led_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => led_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => led_red_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => led_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => led_red_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => led_red_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => led_red_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => led_red_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => led_red_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                  --              (terminated)
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	led_green_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                  --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                      --                    reset.reset
			uav_address              => led_green_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => led_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => led_green_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => led_green_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => led_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => led_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => led_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => led_green_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => led_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => led_green_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => led_green_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => led_green_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => led_green_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => led_green_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	button_pio_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                   --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                       --                    reset.reset
			uav_address              => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => button_pio_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => button_pio_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => button_pio_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => button_pio_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => button_pio_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	switch_pio_s1_translator : component system_0_switch_pio_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                   --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                       --                    reset.reset
			uav_address              => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => switch_pio_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_readdata              => switch_pio_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_write                 => open,                                                                     --              (terminated)
			av_read                  => open,                                                                     --              (terminated)
			av_writedata             => open,                                                                     --              (terminated)
			av_begintransfer         => open,                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                     --              (terminated)
			av_burstcount            => open,                                                                     --              (terminated)
			av_byteenable            => open,                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                     --              (terminated)
			av_lock                  => open,                                                                     --              (terminated)
			av_chipselect            => open,                                                                     --              (terminated)
			av_clken                 => open,                                                                     --              (terminated)
			uav_clken                => '0',                                                                      --              (terminated)
			av_debugaccess           => open,                                                                     --              (terminated)
			av_outputenable          => open,                                                                     --              (terminated)
			uav_response             => open,                                                                     --              (terminated)
			av_response              => "00",                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                       --              (terminated)
		);

	sd_dat_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                   --                    reset.reset
			uav_address              => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sd_dat_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sd_dat_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => sd_dat_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sd_dat_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sd_dat_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	sd_cmd_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                   --                    reset.reset
			uav_address              => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sd_cmd_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sd_cmd_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => sd_cmd_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sd_cmd_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sd_cmd_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	sd_clk_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                               --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                   --                    reset.reset
			uav_address              => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sd_clk_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sd_clk_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => sd_clk_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sd_clk_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => sd_clk_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_byteenable            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			av_clken                 => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	isp1362_hc_translator : component system_0_isp1362_hc_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 3,
			AV_WRITE_WAIT_CYCLES           => 3,
			AV_SETUP_WAIT_CYCLES           => 7,
			AV_DATA_HOLD_CYCLES            => 7
		)
		port map (
			clk                      => clk_50,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                    reset.reset
			uav_address              => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => isp1362_hc_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => isp1362_hc_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => isp1362_hc_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => isp1362_hc_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => isp1362_hc_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => isp1362_hc_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	isp1362_dc_translator : component system_0_isp1362_hc_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 8,
			AV_WRITE_WAIT_CYCLES           => 8,
			AV_SETUP_WAIT_CYCLES           => 8,
			AV_DATA_HOLD_CYCLES            => 8
		)
		port map (
			clk                      => clk_50,                                                                --                      clk.clk
			reset                    => rst_controller_001_reset_out_reset,                                    --                    reset.reset
			uav_address              => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => isp1362_dc_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => isp1362_dc_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => isp1362_dc_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => isp1362_dc_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => isp1362_dc_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => isp1362_dc_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                  --              (terminated)
			av_beginbursttransfer    => open,                                                                  --              (terminated)
			av_burstcount            => open,                                                                  --              (terminated)
			av_byteenable            => open,                                                                  --              (terminated)
			av_readdatavalid         => '0',                                                                   --              (terminated)
			av_waitrequest           => '0',                                                                   --              (terminated)
			av_writebyteenable       => open,                                                                  --              (terminated)
			av_lock                  => open,                                                                  --              (terminated)
			av_clken                 => open,                                                                  --              (terminated)
			uav_clken                => '0',                                                                   --              (terminated)
			av_debugaccess           => open,                                                                  --              (terminated)
			av_outputenable          => open,                                                                  --              (terminated)
			uav_response             => open,                                                                  --              (terminated)
			av_response              => "00",                                                                  --              (terminated)
			uav_writeresponserequest => '0',                                                                   --              (terminated)
			uav_writeresponsevalid   => open,                                                                  --              (terminated)
			av_writeresponserequest  => open,                                                                  --              (terminated)
			av_writeresponsevalid    => '0'                                                                    --              (terminated)
		);

	audio_0_avalon_slave_0_translator : component system_0_audio_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                            --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                --                    reset.reset
			uav_address              => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_write                 => audio_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --      avalon_anti_slave_0.write
			av_readdata              => audio_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => audio_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_address               => open,                                                                              --              (terminated)
			av_read                  => open,                                                                              --              (terminated)
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_byteenable            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_waitrequest           => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_chipselect            => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	vga_0_avalon_slave_0_translator : component system_0_vga_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 19,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 1,
			AV_DATA_HOLD_CYCLES            => 1
		)
		port map (
			clk                      => clk_50,                                                                          --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                              --                    reset.reset
			uav_address              => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => vga_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                            --              (terminated)
			av_beginbursttransfer    => open,                                                                            --              (terminated)
			av_burstcount            => open,                                                                            --              (terminated)
			av_byteenable            => open,                                                                            --              (terminated)
			av_readdatavalid         => '0',                                                                             --              (terminated)
			av_waitrequest           => '0',                                                                             --              (terminated)
			av_writebyteenable       => open,                                                                            --              (terminated)
			av_lock                  => open,                                                                            --              (terminated)
			av_clken                 => open,                                                                            --              (terminated)
			uav_clken                => '0',                                                                             --              (terminated)
			av_debugaccess           => open,                                                                            --              (terminated)
			av_outputenable          => open,                                                                            --              (terminated)
			uav_response             => open,                                                                            --              (terminated)
			av_response              => "00",                                                                            --              (terminated)
			uav_writeresponserequest => '0',                                                                             --              (terminated)
			uav_writeresponsevalid   => open,                                                                            --              (terminated)
			av_writeresponserequest  => open,                                                                            --              (terminated)
			av_writeresponsevalid    => '0'                                                                              --              (terminated)
		);

	dm9000a_avalon_slave_0_translator : component system_0_isp1362_hc_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 2,
			AV_WRITE_WAIT_CYCLES           => 2,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                            --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                --                    reset.reset
			uav_address              => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                              --              (terminated)
			av_beginbursttransfer    => open,                                                                              --              (terminated)
			av_burstcount            => open,                                                                              --              (terminated)
			av_byteenable            => open,                                                                              --              (terminated)
			av_readdatavalid         => '0',                                                                               --              (terminated)
			av_waitrequest           => '0',                                                                               --              (terminated)
			av_writebyteenable       => open,                                                                              --              (terminated)
			av_lock                  => open,                                                                              --              (terminated)
			av_clken                 => open,                                                                              --              (terminated)
			uav_clken                => '0',                                                                               --              (terminated)
			av_debugaccess           => open,                                                                              --              (terminated)
			av_outputenable          => open,                                                                              --              (terminated)
			uav_response             => open,                                                                              --              (terminated)
			av_response              => "00",                                                                              --              (terminated)
			uav_writeresponserequest => '0',                                                                               --              (terminated)
			uav_writeresponsevalid   => open,                                                                              --              (terminated)
			av_writeresponserequest  => open,                                                                              --              (terminated)
			av_writeresponsevalid    => '0'                                                                                --              (terminated)
		);

	seg7_display_avalon_slave_0_translator : component system_0_seg7_display_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                                 --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                     --                    reset.reset
			uav_address              => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_write                 => seg7_display_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --      avalon_anti_slave_0.write
			av_writedata             => seg7_display_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_address               => open,                                                                                   --              (terminated)
			av_read                  => open,                                                                                   --              (terminated)
			av_readdata              => "11011110101011011101111010101101",                                                     --              (terminated)
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_chipselect            => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	sram_0_avalon_slave_0_translator : component system_0_sram_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 18,
			AV_DATA_W                      => 16,
			UAV_DATA_W                     => 16,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 2,
			UAV_BYTEENABLE_W               => 2,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 2,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 2,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 1,
			AV_SETUP_WAIT_CYCLES           => 1,
			AV_DATA_HOLD_CYCLES            => 1
		)
		port map (
			clk                      => clk_50,                                                                           --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                               --                    reset.reset
			uav_address              => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                             --              (terminated)
			av_beginbursttransfer    => open,                                                                             --              (terminated)
			av_burstcount            => open,                                                                             --              (terminated)
			av_readdatavalid         => '0',                                                                              --              (terminated)
			av_waitrequest           => '0',                                                                              --              (terminated)
			av_writebyteenable       => open,                                                                             --              (terminated)
			av_lock                  => open,                                                                             --              (terminated)
			av_clken                 => open,                                                                             --              (terminated)
			uav_clken                => '0',                                                                              --              (terminated)
			av_debugaccess           => open,                                                                             --              (terminated)
			av_outputenable          => open,                                                                             --              (terminated)
			uav_response             => open,                                                                             --              (terminated)
			av_response              => "00",                                                                             --              (terminated)
			uav_writeresponserequest => '0',                                                                              --              (terminated)
			uav_writeresponsevalid   => open,                                                                             --              (terminated)
			av_writeresponserequest  => open,                                                                             --              (terminated)
			av_writeresponsevalid    => '0'                                                                               --              (terminated)
		);

	lab7_final_0_avalon_slave_0_translator : component system_0_lab7_final_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                                 --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                                     --                    reset.reset
			uav_address              => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => lab7_final_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                                   --              (terminated)
			av_burstcount            => open,                                                                                   --              (terminated)
			av_byteenable            => open,                                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                                   --              (terminated)
			av_lock                  => open,                                                                                   --              (terminated)
			av_clken                 => open,                                                                                   --              (terminated)
			uav_clken                => '0',                                                                                    --              (terminated)
			av_debugaccess           => open,                                                                                   --              (terminated)
			av_outputenable          => open,                                                                                   --              (terminated)
			uav_response             => open,                                                                                   --              (terminated)
			av_response              => "00",                                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                                     --              (terminated)
		);

	motor_cw_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                 --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                     --                    reset.reset
			uav_address              => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => motor_cw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => motor_cw_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => motor_cw_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => motor_cw_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => motor_cw_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                   --              (terminated)
			av_begintransfer         => open,                                                                   --              (terminated)
			av_beginbursttransfer    => open,                                                                   --              (terminated)
			av_burstcount            => open,                                                                   --              (terminated)
			av_byteenable            => open,                                                                   --              (terminated)
			av_readdatavalid         => '0',                                                                    --              (terminated)
			av_waitrequest           => '0',                                                                    --              (terminated)
			av_writebyteenable       => open,                                                                   --              (terminated)
			av_lock                  => open,                                                                   --              (terminated)
			av_clken                 => open,                                                                   --              (terminated)
			uav_clken                => '0',                                                                    --              (terminated)
			av_debugaccess           => open,                                                                   --              (terminated)
			av_outputenable          => open,                                                                   --              (terminated)
			uav_response             => open,                                                                   --              (terminated)
			av_response              => "00",                                                                   --              (terminated)
			uav_writeresponserequest => '0',                                                                    --              (terminated)
			uav_writeresponsevalid   => open,                                                                   --              (terminated)
			av_writeresponserequest  => open,                                                                   --              (terminated)
			av_writeresponsevalid    => '0'                                                                     --              (terminated)
		);

	motor_ccw_s1_translator : component system_0_led_red_s1_translator
		generic map (
			AV_ADDRESS_W                   => 2,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 1,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 25,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_50,                                                                  --                      clk.clk
			reset                    => rst_controller_002_reset_out_reset,                                      --                    reset.reset
			uav_address              => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => motor_ccw_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => motor_ccw_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => motor_ccw_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => motor_ccw_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => motor_ccw_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_read                  => open,                                                                    --              (terminated)
			av_begintransfer         => open,                                                                    --              (terminated)
			av_beginbursttransfer    => open,                                                                    --              (terminated)
			av_burstcount            => open,                                                                    --              (terminated)
			av_byteenable            => open,                                                                    --              (terminated)
			av_readdatavalid         => '0',                                                                     --              (terminated)
			av_waitrequest           => '0',                                                                     --              (terminated)
			av_writebyteenable       => open,                                                                    --              (terminated)
			av_lock                  => open,                                                                    --              (terminated)
			av_clken                 => open,                                                                    --              (terminated)
			uav_clken                => '0',                                                                     --              (terminated)
			av_debugaccess           => open,                                                                    --              (terminated)
			av_outputenable          => open,                                                                    --              (terminated)
			uav_response             => open,                                                                    --              (terminated)
			av_response              => "00",                                                                    --              (terminated)
			uav_writeresponserequest => '0',                                                                     --              (terminated)
			uav_writeresponsevalid   => open,                                                                    --              (terminated)
			av_writeresponserequest  => open,                                                                    --              (terminated)
			av_writeresponsevalid    => '0'                                                                      --              (terminated)
		);

	cpu_0_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_THREAD_ID_H           => 92,
			PKT_THREAD_ID_L           => 92,
			PKT_CACHE_H               => 99,
			PKT_CACHE_L               => 96,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			ST_DATA_W                 => 102,
			ST_CHANNEL_W              => 27,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                               --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			av_address              => cpu_0_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_0_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_0_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_0_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_0_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_0_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_0_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_0_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_0_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_0_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_0_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => limiter_rsp_src_valid,                                                                --        rp.valid
			rp_data                 => limiter_rsp_src_data,                                                                 --          .data
			rp_channel              => limiter_rsp_src_channel,                                                              --          .channel
			rp_startofpacket        => limiter_rsp_src_startofpacket,                                                        --          .startofpacket
			rp_endofpacket          => limiter_rsp_src_endofpacket,                                                          --          .endofpacket
			rp_ready                => limiter_rsp_src_ready,                                                                --          .ready
			av_response             => open,                                                                                 -- (terminated)
			av_writeresponserequest => '0',                                                                                  -- (terminated)
			av_writeresponsevalid   => open                                                                                  -- (terminated)
		);

	cpu_0_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_BEGIN_BURST           => 80,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			PKT_BURST_TYPE_H          => 77,
			PKT_BURST_TYPE_L          => 76,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_TRANS_EXCLUSIVE       => 66,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_THREAD_ID_H           => 92,
			PKT_THREAD_ID_L           => 92,
			PKT_CACHE_H               => 99,
			PKT_CACHE_L               => 96,
			PKT_DATA_SIDEBAND_H       => 79,
			PKT_DATA_SIDEBAND_L       => 79,
			PKT_QOS_H                 => 81,
			PKT_QOS_L                 => 81,
			PKT_ADDR_SIDEBAND_H       => 78,
			PKT_ADDR_SIDEBAND_L       => 78,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			ST_DATA_W                 => 102,
			ST_CHANNEL_W              => 27,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 0,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                        --       clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			av_address              => cpu_0_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_0_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_0_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_0_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_0_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_0_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_0_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_0_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_0_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_0_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_0_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                    --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                     --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                  --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                            --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                              --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                    --          .ready
			av_response             => open,                                                                          -- (terminated)
			av_writeresponserequest => '0',                                                                           -- (terminated)
			av_writeresponsevalid   => open                                                                           -- (terminated)
		);

	cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                       --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                           --       clk_reset.reset
			m0_address              => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_src_ready,                                                                       --              cp.ready
			cp_valid                => cmd_xbar_mux_src_valid,                                                                       --                .valid
			cp_data                 => cmd_xbar_mux_src_data,                                                                        --                .data
			cp_startofpacket        => cmd_xbar_mux_src_startofpacket,                                                               --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_src_endofpacket,                                                                 --                .endofpacket
			cp_channel              => cmd_xbar_mux_src_channel,                                                                     --                .channel
			rf_sink_ready           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                         --     (terminated)
			m0_writeresponserequest => open,                                                                                         --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                           --     (terminated)
		);

	cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                       --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                           -- clk_reset.reset
			in_data           => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                         -- (terminated)
			csr_read          => '0',                                                                                          -- (terminated)
			csr_write         => '0',                                                                                          -- (terminated)
			csr_readdata      => open,                                                                                         -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                           -- (terminated)
			almost_full_data  => open,                                                                                         -- (terminated)
			almost_empty_data => open,                                                                                         -- (terminated)
			in_empty          => '0',                                                                                          -- (terminated)
			out_empty         => open,                                                                                         -- (terminated)
			in_error          => '0',                                                                                          -- (terminated)
			out_error         => open,                                                                                         -- (terminated)
			in_channel        => '0',                                                                                          -- (terminated)
			out_channel       => open                                                                                          -- (terminated)
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent : component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 62,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_POSTED          => 44,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			PKT_TRANS_LOCK            => 47,
			PKT_SRC_ID_H              => 68,
			PKT_SRC_ID_L              => 64,
			PKT_DEST_ID_H             => 73,
			PKT_DEST_ID_L             => 69,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_PROTECTION_H          => 77,
			PKT_PROTECTION_L          => 75,
			PKT_RESPONSE_STATUS_H     => 83,
			PKT_RESPONSE_STATUS_L     => 82,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 84,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sdram_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_source0_ready,                                                     --              cp.ready
			cp_valid                => burst_adapter_source0_valid,                                                     --                .valid
			cp_data                 => burst_adapter_source0_data,                                                      --                .data
			cp_startofpacket        => burst_adapter_source0_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => burst_adapter_source0_endofpacket,                                               --                .endofpacket
			cp_channel              => burst_adapter_source0_channel,                                                   --                .channel
			rf_sink_ready           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 85,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sdram_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo : component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 18,
			FIFO_DEPTH          => 8,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 3,
			USE_MEMORY_BLOCKS   => 1,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                    --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                        -- clk_reset.reset
			in_data           => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                      -- (terminated)
			csr_read          => '0',                                                                       -- (terminated)
			csr_write         => '0',                                                                       -- (terminated)
			csr_readdata      => open,                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                        -- (terminated)
			almost_full_data  => open,                                                                      -- (terminated)
			almost_empty_data => open,                                                                      -- (terminated)
			in_startofpacket  => '0',                                                                       -- (terminated)
			in_endofpacket    => '0',                                                                       -- (terminated)
			out_startofpacket => open,                                                                      -- (terminated)
			out_endofpacket   => open,                                                                      -- (terminated)
			in_empty          => '0',                                                                       -- (terminated)
			out_empty         => open,                                                                      -- (terminated)
			in_error          => '0',                                                                       -- (terminated)
			out_error         => open,                                                                      -- (terminated)
			in_channel        => '0',                                                                       -- (terminated)
			out_channel       => open                                                                       -- (terminated)
		);

	epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                                 --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_002_src_ready,                                                                             --              cp.ready
			cp_valid                => cmd_xbar_mux_002_src_valid,                                                                             --                .valid
			cp_data                 => cmd_xbar_mux_002_src_data,                                                                              --                .data
			cp_startofpacket        => cmd_xbar_mux_002_src_startofpacket,                                                                     --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_002_src_endofpacket,                                                                       --                .endofpacket
			cp_channel              => cmd_xbar_mux_002_src_channel,                                                                           --                .channel
			rf_sink_ready           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                                   --     (terminated)
			m0_writeresponserequest => open,                                                                                                   --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                     --     (terminated)
		);

	epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                                 --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                                   -- (terminated)
			csr_read          => '0',                                                                                                    -- (terminated)
			csr_write         => '0',                                                                                                    -- (terminated)
			csr_readdata      => open,                                                                                                   -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                     -- (terminated)
			almost_full_data  => open,                                                                                                   -- (terminated)
			almost_empty_data => open,                                                                                                   -- (terminated)
			in_empty          => '0',                                                                                                    -- (terminated)
			out_empty         => open,                                                                                                   -- (terminated)
			in_error          => '0',                                                                                                    -- (terminated)
			out_error         => open,                                                                                                   -- (terminated)
			in_channel        => '0',                                                                                                    -- (terminated)
			out_channel       => open                                                                                                    -- (terminated)
		);

	cfi_flash_0_uas_translator_avalon_universal_slave_0_agent : component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 7,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 53,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_ADDR_H                => 33,
			PKT_ADDR_L                => 9,
			PKT_TRANS_COMPRESSED_READ => 34,
			PKT_TRANS_POSTED          => 35,
			PKT_TRANS_WRITE           => 36,
			PKT_TRANS_READ            => 37,
			PKT_TRANS_LOCK            => 38,
			PKT_SRC_ID_H              => 59,
			PKT_SRC_ID_L              => 55,
			PKT_DEST_ID_H             => 64,
			PKT_DEST_ID_L             => 60,
			PKT_BURSTWRAP_H           => 45,
			PKT_BURSTWRAP_L           => 43,
			PKT_BYTE_CNT_H            => 42,
			PKT_BYTE_CNT_L            => 40,
			PKT_PROTECTION_H          => 68,
			PKT_PROTECTION_L          => 66,
			PKT_RESPONSE_STATUS_H     => 74,
			PKT_RESPONSE_STATUS_L     => 73,
			PKT_BURST_SIZE_H          => 48,
			PKT_BURST_SIZE_L          => 46,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 75,
			AVS_BURSTCOUNT_W          => 1,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                               --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                   --       clk_reset.reset
			m0_address              => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_001_source0_ready,                                                      --              cp.ready
			cp_valid                => burst_adapter_001_source0_valid,                                                      --                .valid
			cp_data                 => burst_adapter_001_source0_data,                                                       --                .data
			cp_startofpacket        => burst_adapter_001_source0_startofpacket,                                              --                .startofpacket
			cp_endofpacket          => burst_adapter_001_source0_endofpacket,                                                --                .endofpacket
			cp_channel              => burst_adapter_001_source0_channel,                                                    --                .channel
			rf_sink_ready           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid,       --                .valid
			rdata_fifo_sink_data    => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,        --                .data
			rdata_fifo_src_ready    => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                 --     (terminated)
			m0_writeresponserequest => open,                                                                                 --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                   --     (terminated)
		);

	cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 76,
			FIFO_DEPTH          => 4,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                               --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			in_data           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                 -- (terminated)
			csr_read          => '0',                                                                                  -- (terminated)
			csr_write         => '0',                                                                                  -- (terminated)
			csr_readdata      => open,                                                                                 -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                   -- (terminated)
			almost_full_data  => open,                                                                                 -- (terminated)
			almost_empty_data => open,                                                                                 -- (terminated)
			in_empty          => '0',                                                                                  -- (terminated)
			out_empty         => open,                                                                                 -- (terminated)
			in_error          => '0',                                                                                  -- (terminated)
			out_error         => open,                                                                                 -- (terminated)
			in_channel        => '0',                                                                                  -- (terminated)
			out_channel       => open                                                                                  -- (terminated)
		);

	cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo : component system_0_cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 10,
			FIFO_DEPTH          => 4,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 0,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 0,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,  --        in.data
			in_valid          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid, --          .valid
			in_ready          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready, --          .ready
			out_data          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data,  --       out.data
			out_valid         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid, --          .valid
			out_ready         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready, --          .ready
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_startofpacket  => '0',                                                                            -- (terminated)
			in_endofpacket    => '0',                                                                            -- (terminated)
			out_startofpacket => open,                                                                           -- (terminated)
			out_endofpacket   => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                              --       clk_reset.reset
			m0_address              => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_004_src_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_mux_004_src_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_mux_004_src_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_mux_004_src_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_004_src_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_mux_004_src_channel,                                                                    --                .channel
			rf_sink_ready           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                              --     (terminated)
		);

	sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                              -- clk_reset.reset
			in_data           => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                            -- (terminated)
			csr_read          => '0',                                                                                             -- (terminated)
			csr_write         => '0',                                                                                             -- (terminated)
			csr_readdata      => open,                                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                              -- (terminated)
			almost_full_data  => open,                                                                                            -- (terminated)
			almost_empty_data => open,                                                                                            -- (terminated)
			in_empty          => '0',                                                                                             -- (terminated)
			out_empty         => open,                                                                                            -- (terminated)
			in_error          => '0',                                                                                             -- (terminated)
			out_error         => open,                                                                                            -- (terminated)
			in_channel        => '0',                                                                                             -- (terminated)
			out_channel       => open                                                                                             -- (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                                 --       clk_reset.reset
			m0_address              => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src5_ready,                                                                      --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src5_valid,                                                                      --                .valid
			cp_data                 => cmd_xbar_demux_001_src5_data,                                                                       --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src5_startofpacket,                                                              --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src5_endofpacket,                                                                --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src5_channel,                                                                    --                .channel
			rf_sink_ready           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                 --     (terminated)
		);

	jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                                 -- clk_reset.reset
			in_data           => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                 -- (terminated)
			almost_full_data  => open,                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                -- (terminated)
			out_empty         => open,                                                                                               -- (terminated)
			in_error          => '0',                                                                                                -- (terminated)
			out_error         => open,                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                -- (terminated)
			out_channel       => open                                                                                                -- (terminated)
		);

	uart_0_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                         --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => uart_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src6_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src6_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src6_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src6_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src6_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src6_channel,                                                --                .channel
			rf_sink_ready           => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => uart_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => uart_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => uart_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_0_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src7_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src7_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src7_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src7_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src7_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src7_channel,                                                 --                .channel
			rf_sink_ready           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_0_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_0_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => timer_1_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src8_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src8_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src8_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src8_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src8_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src8_channel,                                                 --                .channel
			rf_sink_ready           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => timer_1_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => timer_1_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                         --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                             --       clk_reset.reset
			m0_address              => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src9_ready,                                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src9_valid,                                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src9_data,                                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src9_startofpacket,                                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src9_endofpacket,                                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src9_channel,                                                                --                .channel
			rf_sink_ready           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                             --     (terminated)
		);

	lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                             -- clk_reset.reset
			in_data           => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                           -- (terminated)
			csr_read          => '0',                                                                                            -- (terminated)
			csr_write         => '0',                                                                                            -- (terminated)
			csr_readdata      => open,                                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                             -- (terminated)
			almost_full_data  => open,                                                                                           -- (terminated)
			almost_empty_data => open,                                                                                           -- (terminated)
			in_empty          => '0',                                                                                            -- (terminated)
			out_empty         => open,                                                                                           -- (terminated)
			in_error          => '0',                                                                                            -- (terminated)
			out_error         => open,                                                                                           -- (terminated)
			in_channel        => '0',                                                                                            -- (terminated)
			out_channel       => open                                                                                            -- (terminated)
		);

	led_red_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => led_red_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_red_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_red_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_red_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_red_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_red_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_red_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_red_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_red_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_red_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_red_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_red_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_red_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src10_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src10_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src10_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src10_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src10_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src10_channel,                                                --                .channel
			rf_sink_ready           => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_red_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_red_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_red_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	led_green_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                            --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => led_green_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => led_green_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => led_green_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => led_green_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => led_green_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => led_green_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => led_green_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => led_green_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => led_green_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => led_green_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => led_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => led_green_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => led_green_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => led_green_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => led_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src11_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src11_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src11_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src11_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src11_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src11_channel,                                                  --                .channel
			rf_sink_ready           => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => led_green_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                            --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                -- clk_reset.reset
			in_data           => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => led_green_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => led_green_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	button_pio_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src12_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src12_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_001_src12_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src12_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src12_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src12_channel,                                                   --                .channel
			rf_sink_ready           => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	switch_pio_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                             --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => switch_pio_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src13_ready,                                                     --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src13_valid,                                                     --                .valid
			cp_data                 => cmd_xbar_demux_001_src13_data,                                                      --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src13_startofpacket,                                             --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src13_endofpacket,                                               --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src13_channel,                                                   --                .channel
			rf_sink_ready           => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => switch_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                 --     (terminated)
		);

	switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                             --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => switch_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => switch_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                               -- (terminated)
			csr_read          => '0',                                                                                -- (terminated)
			csr_write         => '0',                                                                                -- (terminated)
			csr_readdata      => open,                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                 -- (terminated)
			almost_full_data  => open,                                                                               -- (terminated)
			almost_empty_data => open,                                                                               -- (terminated)
			in_empty          => '0',                                                                                -- (terminated)
			out_empty         => open,                                                                               -- (terminated)
			in_error          => '0',                                                                                -- (terminated)
			out_error         => open,                                                                               -- (terminated)
			in_channel        => '0',                                                                                -- (terminated)
			out_channel       => open                                                                                -- (terminated)
		);

	sd_dat_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                         --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sd_dat_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src14_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src14_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src14_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src14_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src14_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src14_channel,                                               --                .channel
			rf_sink_ready           => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sd_dat_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sd_dat_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sd_dat_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	sd_cmd_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                         --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sd_cmd_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src15_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src15_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src15_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src15_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src15_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src15_channel,                                               --                .channel
			rf_sink_ready           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	sd_clk_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                         --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                             --       clk_reset.reset
			m0_address              => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sd_clk_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src16_ready,                                                 --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src16_valid,                                                 --                .valid
			cp_data                 => cmd_xbar_demux_001_src16_data,                                                  --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src16_startofpacket,                                         --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src16_endofpacket,                                           --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src16_channel,                                               --                .channel
			rf_sink_ready           => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sd_clk_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                         --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                             -- clk_reset.reset
			in_data           => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sd_clk_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sd_clk_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	isp1362_hc_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => isp1362_hc_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src17_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src17_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src17_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src17_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src17_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src17_channel,                                                --                .channel
			rf_sink_ready           => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => isp1362_hc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => isp1362_hc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => isp1362_hc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	isp1362_dc_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                          --             clk.clk
			reset                   => rst_controller_001_reset_out_reset,                                              --       clk_reset.reset
			m0_address              => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => isp1362_dc_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src18_ready,                                                  --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src18_valid,                                                  --                .valid
			cp_data                 => cmd_xbar_demux_001_src18_data,                                                   --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src18_startofpacket,                                          --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src18_endofpacket,                                            --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src18_channel,                                                --                .channel
			rf_sink_ready           => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => isp1362_dc_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                            --     (terminated)
			m0_writeresponserequest => open,                                                                            --     (terminated)
			m0_writeresponsevalid   => '0'                                                                              --     (terminated)
		);

	isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                          --       clk.clk
			reset             => rst_controller_001_reset_out_reset,                                              -- clk_reset.reset
			in_data           => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => isp1362_dc_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => isp1362_dc_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                            -- (terminated)
			csr_read          => '0',                                                                             -- (terminated)
			csr_write         => '0',                                                                             -- (terminated)
			csr_readdata      => open,                                                                            -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                              -- (terminated)
			almost_full_data  => open,                                                                            -- (terminated)
			almost_empty_data => open,                                                                            -- (terminated)
			in_empty          => '0',                                                                             -- (terminated)
			out_empty         => open,                                                                            -- (terminated)
			in_error          => '0',                                                                             -- (terminated)
			out_error         => open,                                                                            -- (terminated)
			in_channel        => '0',                                                                             -- (terminated)
			out_channel       => open                                                                             -- (terminated)
		);

	audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                      --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src19_ready,                                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src19_valid,                                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src19_data,                                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src19_startofpacket,                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src19_endofpacket,                                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src19_channel,                                                            --                .channel
			rf_sink_ready           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                      --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                    --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                        --       clk_reset.reset
			m0_address              => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src20_ready,                                                            --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src20_valid,                                                            --                .valid
			cp_data                 => cmd_xbar_demux_001_src20_data,                                                             --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src20_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src20_endofpacket,                                                      --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src20_channel,                                                          --                .channel
			rf_sink_ready           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                      --     (terminated)
			m0_writeresponserequest => open,                                                                                      --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                        --     (terminated)
		);

	vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                    --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                        -- clk_reset.reset
			in_data           => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                      -- (terminated)
			csr_read          => '0',                                                                                       -- (terminated)
			csr_write         => '0',                                                                                       -- (terminated)
			csr_readdata      => open,                                                                                      -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                        -- (terminated)
			almost_full_data  => open,                                                                                      -- (terminated)
			almost_empty_data => open,                                                                                      -- (terminated)
			in_empty          => '0',                                                                                       -- (terminated)
			out_empty         => open,                                                                                      -- (terminated)
			in_error          => '0',                                                                                       -- (terminated)
			out_error         => open,                                                                                      -- (terminated)
			in_channel        => '0',                                                                                       -- (terminated)
			out_channel       => open                                                                                       -- (terminated)
		);

	dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                      --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                          --       clk_reset.reset
			m0_address              => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src21_ready,                                                              --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src21_valid,                                                              --                .valid
			cp_data                 => cmd_xbar_demux_001_src21_data,                                                               --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src21_startofpacket,                                                      --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src21_endofpacket,                                                        --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src21_channel,                                                            --                .channel
			rf_sink_ready           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                        --     (terminated)
			m0_writeresponserequest => open,                                                                                        --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                          --     (terminated)
		);

	dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                      --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                          -- clk_reset.reset
			in_data           => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                        -- (terminated)
			csr_read          => '0',                                                                                         -- (terminated)
			csr_write         => '0',                                                                                         -- (terminated)
			csr_readdata      => open,                                                                                        -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                          -- (terminated)
			almost_full_data  => open,                                                                                        -- (terminated)
			almost_empty_data => open,                                                                                        -- (terminated)
			in_empty          => '0',                                                                                         -- (terminated)
			out_empty         => open,                                                                                        -- (terminated)
			in_error          => '0',                                                                                         -- (terminated)
			out_error         => open,                                                                                        -- (terminated)
			in_channel        => '0',                                                                                         -- (terminated)
			out_channel       => open                                                                                         -- (terminated)
		);

	seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                           --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src22_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src22_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src22_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src22_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src22_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src22_channel,                                                                 --                .channel
			rf_sink_ready           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                           --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 15,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 62,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_POSTED          => 44,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			PKT_TRANS_LOCK            => 47,
			PKT_SRC_ID_H              => 68,
			PKT_SRC_ID_L              => 64,
			PKT_DEST_ID_H             => 73,
			PKT_DEST_ID_L             => 69,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_PROTECTION_H          => 77,
			PKT_PROTECTION_L          => 75,
			PKT_RESPONSE_STATUS_H     => 83,
			PKT_RESPONSE_STATUS_L     => 82,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 84,
			AVS_BURSTCOUNT_W          => 2,
			SUPPRESS_0_BYTEEN_CMD     => 1,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                     --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                         --       clk_reset.reset
			m0_address              => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => burst_adapter_002_source0_ready,                                                            --              cp.ready
			cp_valid                => burst_adapter_002_source0_valid,                                                            --                .valid
			cp_data                 => burst_adapter_002_source0_data,                                                             --                .data
			cp_startofpacket        => burst_adapter_002_source0_startofpacket,                                                    --                .startofpacket
			cp_endofpacket          => burst_adapter_002_source0_endofpacket,                                                      --                .endofpacket
			cp_channel              => burst_adapter_002_source0_channel,                                                          --                .channel
			rf_sink_ready           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                       --     (terminated)
			m0_writeresponserequest => open,                                                                                       --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                         --     (terminated)
		);

	sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_sdram_0_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 85,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                     --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                         -- clk_reset.reset
			in_data           => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                       -- (terminated)
			csr_read          => '0',                                                                                        -- (terminated)
			csr_write         => '0',                                                                                        -- (terminated)
			csr_readdata      => open,                                                                                       -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                         -- (terminated)
			almost_full_data  => open,                                                                                       -- (terminated)
			almost_empty_data => open,                                                                                       -- (terminated)
			in_empty          => '0',                                                                                        -- (terminated)
			out_empty         => open,                                                                                       -- (terminated)
			in_error          => '0',                                                                                        -- (terminated)
			out_error         => open,                                                                                       -- (terminated)
			in_channel        => '0',                                                                                        -- (terminated)
			out_channel       => open                                                                                        -- (terminated)
		);

	lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                                           --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                               --       clk_reset.reset
			m0_address              => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src24_ready,                                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src24_valid,                                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src24_data,                                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src24_startofpacket,                                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src24_endofpacket,                                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src24_channel,                                                                 --                .channel
			rf_sink_ready           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                               --     (terminated)
		);

	lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                                           --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                               -- clk_reset.reset
			in_data           => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                             -- (terminated)
			csr_read          => '0',                                                                                              -- (terminated)
			csr_write         => '0',                                                                                              -- (terminated)
			csr_readdata      => open,                                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                               -- (terminated)
			almost_full_data  => open,                                                                                             -- (terminated)
			almost_empty_data => open,                                                                                             -- (terminated)
			in_empty          => '0',                                                                                              -- (terminated)
			out_empty         => open,                                                                                             -- (terminated)
			in_error          => '0',                                                                                              -- (terminated)
			out_error         => open,                                                                                             -- (terminated)
			in_channel        => '0',                                                                                              -- (terminated)
			out_channel       => open                                                                                              -- (terminated)
		);

	motor_cw_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                           --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                               --       clk_reset.reset
			m0_address              => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => motor_cw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src25_ready,                                                   --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src25_valid,                                                   --                .valid
			cp_data                 => cmd_xbar_demux_001_src25_data,                                                    --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src25_startofpacket,                                           --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src25_endofpacket,                                             --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src25_channel,                                                 --                .channel
			rf_sink_ready           => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => motor_cw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                             --     (terminated)
			m0_writeresponserequest => open,                                                                             --     (terminated)
			m0_writeresponsevalid   => '0'                                                                               --     (terminated)
		);

	motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                           --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                               -- clk_reset.reset
			in_data           => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => motor_cw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => motor_cw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                             -- (terminated)
			csr_read          => '0',                                                                              -- (terminated)
			csr_write         => '0',                                                                              -- (terminated)
			csr_readdata      => open,                                                                             -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                               -- (terminated)
			almost_full_data  => open,                                                                             -- (terminated)
			almost_empty_data => open,                                                                             -- (terminated)
			in_empty          => '0',                                                                              -- (terminated)
			out_empty         => open,                                                                             -- (terminated)
			in_error          => '0',                                                                              -- (terminated)
			out_error         => open,                                                                             -- (terminated)
			in_channel        => '0',                                                                              -- (terminated)
			out_channel       => open                                                                              -- (terminated)
		);

	motor_ccw_s1_translator_avalon_universal_slave_0_agent : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 80,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 60,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 61,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			PKT_TRANS_READ            => 64,
			PKT_TRANS_LOCK            => 65,
			PKT_SRC_ID_H              => 86,
			PKT_SRC_ID_L              => 82,
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_BURSTWRAP_H           => 72,
			PKT_BURSTWRAP_L           => 70,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_PROTECTION_H          => 95,
			PKT_PROTECTION_L          => 93,
			PKT_RESPONSE_STATUS_H     => 101,
			PKT_RESPONSE_STATUS_L     => 100,
			PKT_BURST_SIZE_H          => 75,
			PKT_BURST_SIZE_L          => 73,
			ST_CHANNEL_W              => 27,
			ST_DATA_W                 => 102,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_50,                                                                            --             clk.clk
			reset                   => rst_controller_002_reset_out_reset,                                                --       clk_reset.reset
			m0_address              => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => motor_ccw_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_demux_001_src26_ready,                                                    --              cp.ready
			cp_valid                => cmd_xbar_demux_001_src26_valid,                                                    --                .valid
			cp_data                 => cmd_xbar_demux_001_src26_data,                                                     --                .data
			cp_startofpacket        => cmd_xbar_demux_001_src26_startofpacket,                                            --                .startofpacket
			cp_endofpacket          => cmd_xbar_demux_001_src26_endofpacket,                                              --                .endofpacket
			cp_channel              => cmd_xbar_demux_001_src26_channel,                                                  --                .channel
			rf_sink_ready           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                              --     (terminated)
			m0_writeresponserequest => open,                                                                              --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                --     (terminated)
		);

	motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component system_0_cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 103,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_50,                                                                            --       clk.clk
			reset             => rst_controller_002_reset_out_reset,                                                -- clk_reset.reset
			in_data           => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                              -- (terminated)
			csr_read          => '0',                                                                               -- (terminated)
			csr_write         => '0',                                                                               -- (terminated)
			csr_readdata      => open,                                                                              -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                -- (terminated)
			almost_full_data  => open,                                                                              -- (terminated)
			almost_empty_data => open,                                                                              -- (terminated)
			in_empty          => '0',                                                                               -- (terminated)
			out_empty         => open,                                                                              -- (terminated)
			in_error          => '0',                                                                               -- (terminated)
			out_error         => open,                                                                              -- (terminated)
			in_channel        => '0',                                                                               -- (terminated)
			out_channel       => open                                                                               -- (terminated)
		);

	addr_router : component system_0_addr_router
		port map (
			sink_ready         => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_0_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                                --       src.ready
			src_valid          => addr_router_src_valid,                                                                --          .valid
			src_data           => addr_router_src_data,                                                                 --          .data
			src_channel        => addr_router_src_channel,                                                              --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                           --          .endofpacket
		);

	addr_router_001 : component system_0_addr_router_001
		port map (
			sink_ready         => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_0_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                        --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                            -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                     --       src.ready
			src_valid          => addr_router_001_src_valid,                                                     --          .valid
			src_data           => addr_router_001_src_data,                                                      --          .data
			src_channel        => addr_router_001_src_channel,                                                   --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                             --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                                --          .endofpacket
		);

	id_router : component system_0_id_router
		port map (
			sink_ready         => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_0_jtag_debug_module_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                             --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                 -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                                --       src.ready
			src_valid          => id_router_src_valid,                                                                --          .valid
			src_data           => id_router_src_data,                                                                 --          .data
			src_channel        => id_router_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                                           --          .endofpacket
		);

	id_router_001 : component system_0_id_router_001
		port map (
			sink_ready         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sdram_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                               --       src.ready
			src_valid          => id_router_001_src_valid,                                               --          .valid
			src_data           => id_router_001_src_data,                                                --          .data
			src_channel        => id_router_001_src_channel,                                             --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                          --          .endofpacket
		);

	id_router_002 : component system_0_id_router
		port map (
			sink_ready         => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => epcs_controller_epcs_control_port_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                                       --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_002_src_ready,                                                                      --       src.ready
			src_valid          => id_router_002_src_valid,                                                                      --          .valid
			src_data           => id_router_002_src_data,                                                                       --          .data
			src_channel        => id_router_002_src_channel,                                                                    --          .channel
			src_startofpacket  => id_router_002_src_startofpacket,                                                              --          .startofpacket
			src_endofpacket    => id_router_002_src_endofpacket                                                                 --          .endofpacket
		);

	id_router_003 : component system_0_id_router_003
		port map (
			sink_ready         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => cfi_flash_0_uas_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                     --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                         -- clk_reset.reset
			src_ready          => id_router_003_src_ready,                                                    --       src.ready
			src_valid          => id_router_003_src_valid,                                                    --          .valid
			src_data           => id_router_003_src_data,                                                     --          .data
			src_channel        => id_router_003_src_channel,                                                  --          .channel
			src_startofpacket  => id_router_003_src_startofpacket,                                            --          .startofpacket
			src_endofpacket    => id_router_003_src_endofpacket                                               --          .endofpacket
		);

	id_router_004 : component system_0_id_router
		port map (
			sink_ready         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sysid_qsys_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                    -- clk_reset.reset
			src_ready          => id_router_004_src_ready,                                                               --       src.ready
			src_valid          => id_router_004_src_valid,                                                               --          .valid
			src_data           => id_router_004_src_data,                                                                --          .data
			src_channel        => id_router_004_src_channel,                                                             --          .channel
			src_startofpacket  => id_router_004_src_startofpacket,                                                       --          .startofpacket
			src_endofpacket    => id_router_004_src_endofpacket                                                          --          .endofpacket
		);

	id_router_005 : component system_0_id_router_005
		port map (
			sink_ready         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => jtag_uart_0_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                       -- clk_reset.reset
			src_ready          => id_router_005_src_ready,                                                                  --       src.ready
			src_valid          => id_router_005_src_valid,                                                                  --          .valid
			src_data           => id_router_005_src_data,                                                                   --          .data
			src_channel        => id_router_005_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_005_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_005_src_endofpacket                                                             --          .endofpacket
		);

	id_router_006 : component system_0_id_router_005
		port map (
			sink_ready         => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => uart_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_006_src_ready,                                              --       src.ready
			src_valid          => id_router_006_src_valid,                                              --          .valid
			src_data           => id_router_006_src_data,                                               --          .data
			src_channel        => id_router_006_src_channel,                                            --          .channel
			src_startofpacket  => id_router_006_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_006_src_endofpacket                                         --          .endofpacket
		);

	id_router_007 : component system_0_id_router_005
		port map (
			sink_ready         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_0_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_007_src_ready,                                               --       src.ready
			src_valid          => id_router_007_src_valid,                                               --          .valid
			src_data           => id_router_007_src_data,                                                --          .data
			src_channel        => id_router_007_src_channel,                                             --          .channel
			src_startofpacket  => id_router_007_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_007_src_endofpacket                                          --          .endofpacket
		);

	id_router_008 : component system_0_id_router_005
		port map (
			sink_ready         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => timer_1_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_008_src_ready,                                               --       src.ready
			src_valid          => id_router_008_src_valid,                                               --          .valid
			src_data           => id_router_008_src_data,                                                --          .data
			src_channel        => id_router_008_src_channel,                                             --          .channel
			src_startofpacket  => id_router_008_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_008_src_endofpacket                                          --          .endofpacket
		);

	id_router_009 : component system_0_id_router_005
		port map (
			sink_ready         => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lcd_16207_0_control_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                                   -- clk_reset.reset
			src_ready          => id_router_009_src_ready,                                                              --       src.ready
			src_valid          => id_router_009_src_valid,                                                              --          .valid
			src_data           => id_router_009_src_data,                                                               --          .data
			src_channel        => id_router_009_src_channel,                                                            --          .channel
			src_startofpacket  => id_router_009_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => id_router_009_src_endofpacket                                                         --          .endofpacket
		);

	id_router_010 : component system_0_id_router_005
		port map (
			sink_ready         => led_red_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_red_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_red_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_red_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_red_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_010_src_ready,                                               --       src.ready
			src_valid          => id_router_010_src_valid,                                               --          .valid
			src_data           => id_router_010_src_data,                                                --          .data
			src_channel        => id_router_010_src_channel,                                             --          .channel
			src_startofpacket  => id_router_010_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_010_src_endofpacket                                          --          .endofpacket
		);

	id_router_011 : component system_0_id_router_005
		port map (
			sink_ready         => led_green_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => led_green_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => led_green_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => led_green_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => led_green_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                  --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_011_src_ready,                                                 --       src.ready
			src_valid          => id_router_011_src_valid,                                                 --          .valid
			src_data           => id_router_011_src_data,                                                  --          .data
			src_channel        => id_router_011_src_channel,                                               --          .channel
			src_startofpacket  => id_router_011_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_011_src_endofpacket                                            --          .endofpacket
		);

	id_router_012 : component system_0_id_router_005
		port map (
			sink_ready         => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_012_src_ready,                                                  --       src.ready
			src_valid          => id_router_012_src_valid,                                                  --          .valid
			src_data           => id_router_012_src_data,                                                   --          .data
			src_channel        => id_router_012_src_channel,                                                --          .channel
			src_startofpacket  => id_router_012_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_012_src_endofpacket                                             --          .endofpacket
		);

	id_router_013 : component system_0_id_router_005
		port map (
			sink_ready         => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => switch_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                   --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_013_src_ready,                                                  --       src.ready
			src_valid          => id_router_013_src_valid,                                                  --          .valid
			src_data           => id_router_013_src_data,                                                   --          .data
			src_channel        => id_router_013_src_channel,                                                --          .channel
			src_startofpacket  => id_router_013_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_013_src_endofpacket                                             --          .endofpacket
		);

	id_router_014 : component system_0_id_router_005
		port map (
			sink_ready         => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sd_dat_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_014_src_ready,                                              --       src.ready
			src_valid          => id_router_014_src_valid,                                              --          .valid
			src_data           => id_router_014_src_data,                                               --          .data
			src_channel        => id_router_014_src_channel,                                            --          .channel
			src_startofpacket  => id_router_014_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_014_src_endofpacket                                         --          .endofpacket
		);

	id_router_015 : component system_0_id_router_005
		port map (
			sink_ready         => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sd_cmd_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_015_src_ready,                                              --       src.ready
			src_valid          => id_router_015_src_valid,                                              --          .valid
			src_data           => id_router_015_src_data,                                               --          .data
			src_channel        => id_router_015_src_channel,                                            --          .channel
			src_startofpacket  => id_router_015_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_015_src_endofpacket                                         --          .endofpacket
		);

	id_router_016 : component system_0_id_router_005
		port map (
			sink_ready         => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sd_clk_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                               --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                   -- clk_reset.reset
			src_ready          => id_router_016_src_ready,                                              --       src.ready
			src_valid          => id_router_016_src_valid,                                              --          .valid
			src_data           => id_router_016_src_data,                                               --          .data
			src_channel        => id_router_016_src_channel,                                            --          .channel
			src_startofpacket  => id_router_016_src_startofpacket,                                      --          .startofpacket
			src_endofpacket    => id_router_016_src_endofpacket                                         --          .endofpacket
		);

	id_router_017 : component system_0_id_router_005
		port map (
			sink_ready         => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => isp1362_hc_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_017_src_ready,                                               --       src.ready
			src_valid          => id_router_017_src_valid,                                               --          .valid
			src_data           => id_router_017_src_data,                                                --          .data
			src_channel        => id_router_017_src_channel,                                             --          .channel
			src_startofpacket  => id_router_017_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_017_src_endofpacket                                          --          .endofpacket
		);

	id_router_018 : component system_0_id_router_005
		port map (
			sink_ready         => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => isp1362_dc_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,                                    -- clk_reset.reset
			src_ready          => id_router_018_src_ready,                                               --       src.ready
			src_valid          => id_router_018_src_valid,                                               --          .valid
			src_data           => id_router_018_src_data,                                                --          .data
			src_channel        => id_router_018_src_channel,                                             --          .channel
			src_startofpacket  => id_router_018_src_startofpacket,                                       --          .startofpacket
			src_endofpacket    => id_router_018_src_endofpacket                                          --          .endofpacket
		);

	id_router_019 : component system_0_id_router_005
		port map (
			sink_ready         => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => audio_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                            --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_019_src_ready,                                                           --       src.ready
			src_valid          => id_router_019_src_valid,                                                           --          .valid
			src_data           => id_router_019_src_data,                                                            --          .data
			src_channel        => id_router_019_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_019_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_019_src_endofpacket                                                      --          .endofpacket
		);

	id_router_020 : component system_0_id_router_005
		port map (
			sink_ready         => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => vga_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                          --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => id_router_020_src_ready,                                                         --       src.ready
			src_valid          => id_router_020_src_valid,                                                         --          .valid
			src_data           => id_router_020_src_data,                                                          --          .data
			src_channel        => id_router_020_src_channel,                                                       --          .channel
			src_startofpacket  => id_router_020_src_startofpacket,                                                 --          .startofpacket
			src_endofpacket    => id_router_020_src_endofpacket                                                    --          .endofpacket
		);

	id_router_021 : component system_0_id_router_005
		port map (
			sink_ready         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => dm9000a_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                            --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                -- clk_reset.reset
			src_ready          => id_router_021_src_ready,                                                           --       src.ready
			src_valid          => id_router_021_src_valid,                                                           --          .valid
			src_data           => id_router_021_src_data,                                                            --          .data
			src_channel        => id_router_021_src_channel,                                                         --          .channel
			src_startofpacket  => id_router_021_src_startofpacket,                                                   --          .startofpacket
			src_endofpacket    => id_router_021_src_endofpacket                                                      --          .endofpacket
		);

	id_router_022 : component system_0_id_router_005
		port map (
			sink_ready         => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => seg7_display_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                                 --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_022_src_ready,                                                                --       src.ready
			src_valid          => id_router_022_src_valid,                                                                --          .valid
			src_data           => id_router_022_src_data,                                                                 --          .data
			src_channel        => id_router_022_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_022_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_022_src_endofpacket                                                           --          .endofpacket
		);

	id_router_023 : component system_0_id_router_023
		port map (
			sink_ready         => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => sram_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                           --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                               -- clk_reset.reset
			src_ready          => id_router_023_src_ready,                                                          --       src.ready
			src_valid          => id_router_023_src_valid,                                                          --          .valid
			src_data           => id_router_023_src_data,                                                           --          .data
			src_channel        => id_router_023_src_channel,                                                        --          .channel
			src_startofpacket  => id_router_023_src_startofpacket,                                                  --          .startofpacket
			src_endofpacket    => id_router_023_src_endofpacket                                                     --          .endofpacket
		);

	id_router_024 : component system_0_id_router_005
		port map (
			sink_ready         => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => lab7_final_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                                 --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => id_router_024_src_ready,                                                                --       src.ready
			src_valid          => id_router_024_src_valid,                                                                --          .valid
			src_data           => id_router_024_src_data,                                                                 --          .data
			src_channel        => id_router_024_src_channel,                                                              --          .channel
			src_startofpacket  => id_router_024_src_startofpacket,                                                        --          .startofpacket
			src_endofpacket    => id_router_024_src_endofpacket                                                           --          .endofpacket
		);

	id_router_025 : component system_0_id_router_005
		port map (
			sink_ready         => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => motor_cw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                 --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                     -- clk_reset.reset
			src_ready          => id_router_025_src_ready,                                                --       src.ready
			src_valid          => id_router_025_src_valid,                                                --          .valid
			src_data           => id_router_025_src_data,                                                 --          .data
			src_channel        => id_router_025_src_channel,                                              --          .channel
			src_startofpacket  => id_router_025_src_startofpacket,                                        --          .startofpacket
			src_endofpacket    => id_router_025_src_endofpacket                                           --          .endofpacket
		);

	id_router_026 : component system_0_id_router_005
		port map (
			sink_ready         => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => motor_ccw_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_50,                                                                  --       clk.clk
			reset              => rst_controller_002_reset_out_reset,                                      -- clk_reset.reset
			src_ready          => id_router_026_src_ready,                                                 --       src.ready
			src_valid          => id_router_026_src_valid,                                                 --          .valid
			src_data           => id_router_026_src_data,                                                  --          .data
			src_channel        => id_router_026_src_channel,                                               --          .channel
			src_startofpacket  => id_router_026_src_startofpacket,                                         --          .startofpacket
			src_endofpacket    => id_router_026_src_endofpacket                                            --          .endofpacket
		);

	limiter : component altera_merlin_traffic_limiter
		generic map (
			PKT_DEST_ID_H             => 91,
			PKT_DEST_ID_L             => 87,
			PKT_TRANS_POSTED          => 62,
			PKT_TRANS_WRITE           => 63,
			MAX_OUTSTANDING_RESPONSES => 9,
			PIPELINED                 => 0,
			ST_DATA_W                 => 102,
			ST_CHANNEL_W              => 27,
			VALID_WIDTH               => 27,
			ENFORCE_ORDER             => 1,
			PREVENT_HAZARDS           => 0,
			PKT_BYTE_CNT_H            => 69,
			PKT_BYTE_CNT_L            => 67,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32
		)
		port map (
			clk                    => clk_50,                             --       clk.clk
			reset                  => rst_controller_001_reset_out_reset, -- clk_reset.reset
			cmd_sink_ready         => addr_router_src_ready,              --  cmd_sink.ready
			cmd_sink_valid         => addr_router_src_valid,              --          .valid
			cmd_sink_data          => addr_router_src_data,               --          .data
			cmd_sink_channel       => addr_router_src_channel,            --          .channel
			cmd_sink_startofpacket => addr_router_src_startofpacket,      --          .startofpacket
			cmd_sink_endofpacket   => addr_router_src_endofpacket,        --          .endofpacket
			cmd_src_ready          => limiter_cmd_src_ready,              --   cmd_src.ready
			cmd_src_data           => limiter_cmd_src_data,               --          .data
			cmd_src_channel        => limiter_cmd_src_channel,            --          .channel
			cmd_src_startofpacket  => limiter_cmd_src_startofpacket,      --          .startofpacket
			cmd_src_endofpacket    => limiter_cmd_src_endofpacket,        --          .endofpacket
			rsp_sink_ready         => rsp_xbar_mux_src_ready,             --  rsp_sink.ready
			rsp_sink_valid         => rsp_xbar_mux_src_valid,             --          .valid
			rsp_sink_channel       => rsp_xbar_mux_src_channel,           --          .channel
			rsp_sink_data          => rsp_xbar_mux_src_data,              --          .data
			rsp_sink_startofpacket => rsp_xbar_mux_src_startofpacket,     --          .startofpacket
			rsp_sink_endofpacket   => rsp_xbar_mux_src_endofpacket,       --          .endofpacket
			rsp_src_ready          => limiter_rsp_src_ready,              --   rsp_src.ready
			rsp_src_valid          => limiter_rsp_src_valid,              --          .valid
			rsp_src_data           => limiter_rsp_src_data,               --          .data
			rsp_src_channel        => limiter_rsp_src_channel,            --          .channel
			rsp_src_startofpacket  => limiter_rsp_src_startofpacket,      --          .startofpacket
			rsp_src_endofpacket    => limiter_rsp_src_endofpacket,        --          .endofpacket
			cmd_src_valid          => limiter_cmd_valid_data              -- cmd_valid.data
		);

	burst_adapter : component system_0_burst_adapter
		generic map (
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 62,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			PKT_BURST_TYPE_H          => 59,
			PKT_BURST_TYPE_L          => 58,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 84,
			ST_CHANNEL_W              => 27,
			OUT_BYTE_CNT_H            => 50,
			OUT_BURSTWRAP_H           => 54,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => clk_50,                              --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,  -- cr0_reset.reset
			sink0_valid           => width_adapter_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_src_data,              --          .data
			sink0_channel         => width_adapter_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_src_ready,             --          .ready
			source0_valid         => burst_adapter_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_source0_data,          --          .data
			source0_channel       => burst_adapter_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_source0_ready          --          .ready
		);

	burst_adapter_001 : component system_0_burst_adapter_001
		generic map (
			PKT_ADDR_H                => 33,
			PKT_ADDR_L                => 9,
			PKT_BEGIN_BURST           => 53,
			PKT_BYTE_CNT_H            => 42,
			PKT_BYTE_CNT_L            => 40,
			PKT_BYTEEN_H              => 8,
			PKT_BYTEEN_L              => 8,
			PKT_BURST_SIZE_H          => 48,
			PKT_BURST_SIZE_L          => 46,
			PKT_BURST_TYPE_H          => 50,
			PKT_BURST_TYPE_L          => 49,
			PKT_BURSTWRAP_H           => 45,
			PKT_BURSTWRAP_L           => 43,
			PKT_TRANS_COMPRESSED_READ => 34,
			PKT_TRANS_WRITE           => 36,
			PKT_TRANS_READ            => 37,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 75,
			ST_CHANNEL_W              => 27,
			OUT_BYTE_CNT_H            => 40,
			OUT_BURSTWRAP_H           => 45,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 3,
			BURSTWRAP_CONST_VALUE     => 3
		)
		port map (
			clk                   => clk_50,                                  --       cr0.clk
			reset                 => rst_controller_001_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_002_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_002_src_data,              --          .data
			sink0_channel         => width_adapter_002_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_002_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_002_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_002_src_ready,             --          .ready
			source0_valid         => burst_adapter_001_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_001_source0_data,          --          .data
			source0_channel       => burst_adapter_001_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_001_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_001_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_001_source0_ready          --          .ready
		);

	burst_adapter_002 : component system_0_burst_adapter
		generic map (
			PKT_ADDR_H                => 42,
			PKT_ADDR_L                => 18,
			PKT_BEGIN_BURST           => 62,
			PKT_BYTE_CNT_H            => 51,
			PKT_BYTE_CNT_L            => 49,
			PKT_BYTEEN_H              => 17,
			PKT_BYTEEN_L              => 16,
			PKT_BURST_SIZE_H          => 57,
			PKT_BURST_SIZE_L          => 55,
			PKT_BURST_TYPE_H          => 59,
			PKT_BURST_TYPE_L          => 58,
			PKT_BURSTWRAP_H           => 54,
			PKT_BURSTWRAP_L           => 52,
			PKT_TRANS_COMPRESSED_READ => 43,
			PKT_TRANS_WRITE           => 45,
			PKT_TRANS_READ            => 46,
			OUT_NARROW_SIZE           => 0,
			IN_NARROW_SIZE            => 0,
			OUT_FIXED                 => 0,
			OUT_COMPLETE_WRAP         => 0,
			ST_DATA_W                 => 84,
			ST_CHANNEL_W              => 27,
			OUT_BYTE_CNT_H            => 50,
			OUT_BURSTWRAP_H           => 54,
			COMPRESSED_READ_SUPPORT   => 0,
			BYTEENABLE_SYNTHESIS      => 1,
			PIPE_INPUTS               => 0,
			NO_WRAP_SUPPORT           => 0,
			BURSTWRAP_CONST_MASK      => 7,
			BURSTWRAP_CONST_VALUE     => 7
		)
		port map (
			clk                   => clk_50,                                  --       cr0.clk
			reset                 => rst_controller_002_reset_out_reset,      -- cr0_reset.reset
			sink0_valid           => width_adapter_004_src_valid,             --     sink0.valid
			sink0_data            => width_adapter_004_src_data,              --          .data
			sink0_channel         => width_adapter_004_src_channel,           --          .channel
			sink0_startofpacket   => width_adapter_004_src_startofpacket,     --          .startofpacket
			sink0_endofpacket     => width_adapter_004_src_endofpacket,       --          .endofpacket
			sink0_ready           => width_adapter_004_src_ready,             --          .ready
			source0_valid         => burst_adapter_002_source0_valid,         --   source0.valid
			source0_data          => burst_adapter_002_source0_data,          --          .data
			source0_channel       => burst_adapter_002_source0_channel,       --          .channel
			source0_startofpacket => burst_adapter_002_source0_startofpacket, --          .startofpacket
			source0_endofpacket   => burst_adapter_002_source0_endofpacket,   --          .endofpacket
			source0_ready         => burst_adapter_002_source0_ready          --          .ready
		);

	rst_controller : component system_0_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "none",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                   -- reset_in0.reset
			reset_in1  => cpu_0_jtag_debug_module_reset_reset, -- reset_in1.reset
			clk        => open,                                --       clk.clk
			reset_out  => open,                                -- reset_out.reset
			reset_req  => open,                                -- (terminated)
			reset_in2  => '0',                                 -- (terminated)
			reset_in3  => '0',                                 -- (terminated)
			reset_in4  => '0',                                 -- (terminated)
			reset_in5  => '0',                                 -- (terminated)
			reset_in6  => '0',                                 -- (terminated)
			reset_in7  => '0',                                 -- (terminated)
			reset_in8  => '0',                                 -- (terminated)
			reset_in9  => '0',                                 -- (terminated)
			reset_in10 => '0',                                 -- (terminated)
			reset_in11 => '0',                                 -- (terminated)
			reset_in12 => '0',                                 -- (terminated)
			reset_in13 => '0',                                 -- (terminated)
			reset_in14 => '0',                                 -- (terminated)
			reset_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component system_0_rst_controller
		generic map (
			NUM_RESET_INPUTS        => 2,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => cpu_0_jtag_debug_module_reset_reset, -- reset_in0.reset
			reset_in1  => reset_n_ports_inv,                   -- reset_in1.reset
			clk        => clk_50,                              --       clk.clk
			reset_out  => rst_controller_001_reset_out_reset,  -- reset_out.reset
			reset_req  => open,                                -- (terminated)
			reset_in2  => '0',                                 -- (terminated)
			reset_in3  => '0',                                 -- (terminated)
			reset_in4  => '0',                                 -- (terminated)
			reset_in5  => '0',                                 -- (terminated)
			reset_in6  => '0',                                 -- (terminated)
			reset_in7  => '0',                                 -- (terminated)
			reset_in8  => '0',                                 -- (terminated)
			reset_in9  => '0',                                 -- (terminated)
			reset_in10 => '0',                                 -- (terminated)
			reset_in11 => '0',                                 -- (terminated)
			reset_in12 => '0',                                 -- (terminated)
			reset_in13 => '0',                                 -- (terminated)
			reset_in14 => '0',                                 -- (terminated)
			reset_in15 => '0'                                  -- (terminated)
		);

	rst_controller_002 : component system_0_rst_controller_002
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 0
		)
		port map (
			reset_in0  => reset_n_ports_inv,                  -- reset_in0.reset
			clk        => clk_50,                             --       clk.clk
			reset_out  => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req  => open,                               -- (terminated)
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component system_0_cmd_xbar_demux
		port map (
			clk                => clk_50,                             --        clk.clk
			reset              => rst_controller_001_reset_out_reset, --  clk_reset.reset
			sink_ready         => limiter_cmd_src_ready,              --       sink.ready
			sink_channel       => limiter_cmd_src_channel,            --           .channel
			sink_data          => limiter_cmd_src_data,               --           .data
			sink_startofpacket => limiter_cmd_src_startofpacket,      --           .startofpacket
			sink_endofpacket   => limiter_cmd_src_endofpacket,        --           .endofpacket
			sink_valid         => limiter_cmd_valid_data,             -- sink_valid.data
			src0_ready         => cmd_xbar_demux_src0_ready,          --       src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,          --           .valid
			src0_data          => cmd_xbar_demux_src0_data,           --           .data
			src0_channel       => cmd_xbar_demux_src0_channel,        --           .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket,  --           .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,    --           .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,          --       src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,          --           .valid
			src1_data          => cmd_xbar_demux_src1_data,           --           .data
			src1_channel       => cmd_xbar_demux_src1_channel,        --           .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket,  --           .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket,    --           .endofpacket
			src2_ready         => cmd_xbar_demux_src2_ready,          --       src2.ready
			src2_valid         => cmd_xbar_demux_src2_valid,          --           .valid
			src2_data          => cmd_xbar_demux_src2_data,           --           .data
			src2_channel       => cmd_xbar_demux_src2_channel,        --           .channel
			src2_startofpacket => cmd_xbar_demux_src2_startofpacket,  --           .startofpacket
			src2_endofpacket   => cmd_xbar_demux_src2_endofpacket,    --           .endofpacket
			src3_ready         => cmd_xbar_demux_src3_ready,          --       src3.ready
			src3_valid         => cmd_xbar_demux_src3_valid,          --           .valid
			src3_data          => cmd_xbar_demux_src3_data,           --           .data
			src3_channel       => cmd_xbar_demux_src3_channel,        --           .channel
			src3_startofpacket => cmd_xbar_demux_src3_startofpacket,  --           .startofpacket
			src3_endofpacket   => cmd_xbar_demux_src3_endofpacket,    --           .endofpacket
			src4_ready         => cmd_xbar_demux_src4_ready,          --       src4.ready
			src4_valid         => cmd_xbar_demux_src4_valid,          --           .valid
			src4_data          => cmd_xbar_demux_src4_data,           --           .data
			src4_channel       => cmd_xbar_demux_src4_channel,        --           .channel
			src4_startofpacket => cmd_xbar_demux_src4_startofpacket,  --           .startofpacket
			src4_endofpacket   => cmd_xbar_demux_src4_endofpacket     --           .endofpacket
		);

	cmd_xbar_demux_001 : component system_0_cmd_xbar_demux_001
		port map (
			clk                 => clk_50,                                 --       clk.clk
			reset               => rst_controller_001_reset_out_reset,     -- clk_reset.reset
			sink_ready          => addr_router_001_src_ready,              --      sink.ready
			sink_channel        => addr_router_001_src_channel,            --          .channel
			sink_data           => addr_router_001_src_data,               --          .data
			sink_startofpacket  => addr_router_001_src_startofpacket,      --          .startofpacket
			sink_endofpacket    => addr_router_001_src_endofpacket,        --          .endofpacket
			sink_valid(0)       => addr_router_001_src_valid,              --          .valid
			src0_ready          => cmd_xbar_demux_001_src0_ready,          --      src0.ready
			src0_valid          => cmd_xbar_demux_001_src0_valid,          --          .valid
			src0_data           => cmd_xbar_demux_001_src0_data,           --          .data
			src0_channel        => cmd_xbar_demux_001_src0_channel,        --          .channel
			src0_startofpacket  => cmd_xbar_demux_001_src0_startofpacket,  --          .startofpacket
			src0_endofpacket    => cmd_xbar_demux_001_src0_endofpacket,    --          .endofpacket
			src1_ready          => cmd_xbar_demux_001_src1_ready,          --      src1.ready
			src1_valid          => cmd_xbar_demux_001_src1_valid,          --          .valid
			src1_data           => cmd_xbar_demux_001_src1_data,           --          .data
			src1_channel        => cmd_xbar_demux_001_src1_channel,        --          .channel
			src1_startofpacket  => cmd_xbar_demux_001_src1_startofpacket,  --          .startofpacket
			src1_endofpacket    => cmd_xbar_demux_001_src1_endofpacket,    --          .endofpacket
			src2_ready          => cmd_xbar_demux_001_src2_ready,          --      src2.ready
			src2_valid          => cmd_xbar_demux_001_src2_valid,          --          .valid
			src2_data           => cmd_xbar_demux_001_src2_data,           --          .data
			src2_channel        => cmd_xbar_demux_001_src2_channel,        --          .channel
			src2_startofpacket  => cmd_xbar_demux_001_src2_startofpacket,  --          .startofpacket
			src2_endofpacket    => cmd_xbar_demux_001_src2_endofpacket,    --          .endofpacket
			src3_ready          => cmd_xbar_demux_001_src3_ready,          --      src3.ready
			src3_valid          => cmd_xbar_demux_001_src3_valid,          --          .valid
			src3_data           => cmd_xbar_demux_001_src3_data,           --          .data
			src3_channel        => cmd_xbar_demux_001_src3_channel,        --          .channel
			src3_startofpacket  => cmd_xbar_demux_001_src3_startofpacket,  --          .startofpacket
			src3_endofpacket    => cmd_xbar_demux_001_src3_endofpacket,    --          .endofpacket
			src4_ready          => cmd_xbar_demux_001_src4_ready,          --      src4.ready
			src4_valid          => cmd_xbar_demux_001_src4_valid,          --          .valid
			src4_data           => cmd_xbar_demux_001_src4_data,           --          .data
			src4_channel        => cmd_xbar_demux_001_src4_channel,        --          .channel
			src4_startofpacket  => cmd_xbar_demux_001_src4_startofpacket,  --          .startofpacket
			src4_endofpacket    => cmd_xbar_demux_001_src4_endofpacket,    --          .endofpacket
			src5_ready          => cmd_xbar_demux_001_src5_ready,          --      src5.ready
			src5_valid          => cmd_xbar_demux_001_src5_valid,          --          .valid
			src5_data           => cmd_xbar_demux_001_src5_data,           --          .data
			src5_channel        => cmd_xbar_demux_001_src5_channel,        --          .channel
			src5_startofpacket  => cmd_xbar_demux_001_src5_startofpacket,  --          .startofpacket
			src5_endofpacket    => cmd_xbar_demux_001_src5_endofpacket,    --          .endofpacket
			src6_ready          => cmd_xbar_demux_001_src6_ready,          --      src6.ready
			src6_valid          => cmd_xbar_demux_001_src6_valid,          --          .valid
			src6_data           => cmd_xbar_demux_001_src6_data,           --          .data
			src6_channel        => cmd_xbar_demux_001_src6_channel,        --          .channel
			src6_startofpacket  => cmd_xbar_demux_001_src6_startofpacket,  --          .startofpacket
			src6_endofpacket    => cmd_xbar_demux_001_src6_endofpacket,    --          .endofpacket
			src7_ready          => cmd_xbar_demux_001_src7_ready,          --      src7.ready
			src7_valid          => cmd_xbar_demux_001_src7_valid,          --          .valid
			src7_data           => cmd_xbar_demux_001_src7_data,           --          .data
			src7_channel        => cmd_xbar_demux_001_src7_channel,        --          .channel
			src7_startofpacket  => cmd_xbar_demux_001_src7_startofpacket,  --          .startofpacket
			src7_endofpacket    => cmd_xbar_demux_001_src7_endofpacket,    --          .endofpacket
			src8_ready          => cmd_xbar_demux_001_src8_ready,          --      src8.ready
			src8_valid          => cmd_xbar_demux_001_src8_valid,          --          .valid
			src8_data           => cmd_xbar_demux_001_src8_data,           --          .data
			src8_channel        => cmd_xbar_demux_001_src8_channel,        --          .channel
			src8_startofpacket  => cmd_xbar_demux_001_src8_startofpacket,  --          .startofpacket
			src8_endofpacket    => cmd_xbar_demux_001_src8_endofpacket,    --          .endofpacket
			src9_ready          => cmd_xbar_demux_001_src9_ready,          --      src9.ready
			src9_valid          => cmd_xbar_demux_001_src9_valid,          --          .valid
			src9_data           => cmd_xbar_demux_001_src9_data,           --          .data
			src9_channel        => cmd_xbar_demux_001_src9_channel,        --          .channel
			src9_startofpacket  => cmd_xbar_demux_001_src9_startofpacket,  --          .startofpacket
			src9_endofpacket    => cmd_xbar_demux_001_src9_endofpacket,    --          .endofpacket
			src10_ready         => cmd_xbar_demux_001_src10_ready,         --     src10.ready
			src10_valid         => cmd_xbar_demux_001_src10_valid,         --          .valid
			src10_data          => cmd_xbar_demux_001_src10_data,          --          .data
			src10_channel       => cmd_xbar_demux_001_src10_channel,       --          .channel
			src10_startofpacket => cmd_xbar_demux_001_src10_startofpacket, --          .startofpacket
			src10_endofpacket   => cmd_xbar_demux_001_src10_endofpacket,   --          .endofpacket
			src11_ready         => cmd_xbar_demux_001_src11_ready,         --     src11.ready
			src11_valid         => cmd_xbar_demux_001_src11_valid,         --          .valid
			src11_data          => cmd_xbar_demux_001_src11_data,          --          .data
			src11_channel       => cmd_xbar_demux_001_src11_channel,       --          .channel
			src11_startofpacket => cmd_xbar_demux_001_src11_startofpacket, --          .startofpacket
			src11_endofpacket   => cmd_xbar_demux_001_src11_endofpacket,   --          .endofpacket
			src12_ready         => cmd_xbar_demux_001_src12_ready,         --     src12.ready
			src12_valid         => cmd_xbar_demux_001_src12_valid,         --          .valid
			src12_data          => cmd_xbar_demux_001_src12_data,          --          .data
			src12_channel       => cmd_xbar_demux_001_src12_channel,       --          .channel
			src12_startofpacket => cmd_xbar_demux_001_src12_startofpacket, --          .startofpacket
			src12_endofpacket   => cmd_xbar_demux_001_src12_endofpacket,   --          .endofpacket
			src13_ready         => cmd_xbar_demux_001_src13_ready,         --     src13.ready
			src13_valid         => cmd_xbar_demux_001_src13_valid,         --          .valid
			src13_data          => cmd_xbar_demux_001_src13_data,          --          .data
			src13_channel       => cmd_xbar_demux_001_src13_channel,       --          .channel
			src13_startofpacket => cmd_xbar_demux_001_src13_startofpacket, --          .startofpacket
			src13_endofpacket   => cmd_xbar_demux_001_src13_endofpacket,   --          .endofpacket
			src14_ready         => cmd_xbar_demux_001_src14_ready,         --     src14.ready
			src14_valid         => cmd_xbar_demux_001_src14_valid,         --          .valid
			src14_data          => cmd_xbar_demux_001_src14_data,          --          .data
			src14_channel       => cmd_xbar_demux_001_src14_channel,       --          .channel
			src14_startofpacket => cmd_xbar_demux_001_src14_startofpacket, --          .startofpacket
			src14_endofpacket   => cmd_xbar_demux_001_src14_endofpacket,   --          .endofpacket
			src15_ready         => cmd_xbar_demux_001_src15_ready,         --     src15.ready
			src15_valid         => cmd_xbar_demux_001_src15_valid,         --          .valid
			src15_data          => cmd_xbar_demux_001_src15_data,          --          .data
			src15_channel       => cmd_xbar_demux_001_src15_channel,       --          .channel
			src15_startofpacket => cmd_xbar_demux_001_src15_startofpacket, --          .startofpacket
			src15_endofpacket   => cmd_xbar_demux_001_src15_endofpacket,   --          .endofpacket
			src16_ready         => cmd_xbar_demux_001_src16_ready,         --     src16.ready
			src16_valid         => cmd_xbar_demux_001_src16_valid,         --          .valid
			src16_data          => cmd_xbar_demux_001_src16_data,          --          .data
			src16_channel       => cmd_xbar_demux_001_src16_channel,       --          .channel
			src16_startofpacket => cmd_xbar_demux_001_src16_startofpacket, --          .startofpacket
			src16_endofpacket   => cmd_xbar_demux_001_src16_endofpacket,   --          .endofpacket
			src17_ready         => cmd_xbar_demux_001_src17_ready,         --     src17.ready
			src17_valid         => cmd_xbar_demux_001_src17_valid,         --          .valid
			src17_data          => cmd_xbar_demux_001_src17_data,          --          .data
			src17_channel       => cmd_xbar_demux_001_src17_channel,       --          .channel
			src17_startofpacket => cmd_xbar_demux_001_src17_startofpacket, --          .startofpacket
			src17_endofpacket   => cmd_xbar_demux_001_src17_endofpacket,   --          .endofpacket
			src18_ready         => cmd_xbar_demux_001_src18_ready,         --     src18.ready
			src18_valid         => cmd_xbar_demux_001_src18_valid,         --          .valid
			src18_data          => cmd_xbar_demux_001_src18_data,          --          .data
			src18_channel       => cmd_xbar_demux_001_src18_channel,       --          .channel
			src18_startofpacket => cmd_xbar_demux_001_src18_startofpacket, --          .startofpacket
			src18_endofpacket   => cmd_xbar_demux_001_src18_endofpacket,   --          .endofpacket
			src19_ready         => cmd_xbar_demux_001_src19_ready,         --     src19.ready
			src19_valid         => cmd_xbar_demux_001_src19_valid,         --          .valid
			src19_data          => cmd_xbar_demux_001_src19_data,          --          .data
			src19_channel       => cmd_xbar_demux_001_src19_channel,       --          .channel
			src19_startofpacket => cmd_xbar_demux_001_src19_startofpacket, --          .startofpacket
			src19_endofpacket   => cmd_xbar_demux_001_src19_endofpacket,   --          .endofpacket
			src20_ready         => cmd_xbar_demux_001_src20_ready,         --     src20.ready
			src20_valid         => cmd_xbar_demux_001_src20_valid,         --          .valid
			src20_data          => cmd_xbar_demux_001_src20_data,          --          .data
			src20_channel       => cmd_xbar_demux_001_src20_channel,       --          .channel
			src20_startofpacket => cmd_xbar_demux_001_src20_startofpacket, --          .startofpacket
			src20_endofpacket   => cmd_xbar_demux_001_src20_endofpacket,   --          .endofpacket
			src21_ready         => cmd_xbar_demux_001_src21_ready,         --     src21.ready
			src21_valid         => cmd_xbar_demux_001_src21_valid,         --          .valid
			src21_data          => cmd_xbar_demux_001_src21_data,          --          .data
			src21_channel       => cmd_xbar_demux_001_src21_channel,       --          .channel
			src21_startofpacket => cmd_xbar_demux_001_src21_startofpacket, --          .startofpacket
			src21_endofpacket   => cmd_xbar_demux_001_src21_endofpacket,   --          .endofpacket
			src22_ready         => cmd_xbar_demux_001_src22_ready,         --     src22.ready
			src22_valid         => cmd_xbar_demux_001_src22_valid,         --          .valid
			src22_data          => cmd_xbar_demux_001_src22_data,          --          .data
			src22_channel       => cmd_xbar_demux_001_src22_channel,       --          .channel
			src22_startofpacket => cmd_xbar_demux_001_src22_startofpacket, --          .startofpacket
			src22_endofpacket   => cmd_xbar_demux_001_src22_endofpacket,   --          .endofpacket
			src23_ready         => cmd_xbar_demux_001_src23_ready,         --     src23.ready
			src23_valid         => cmd_xbar_demux_001_src23_valid,         --          .valid
			src23_data          => cmd_xbar_demux_001_src23_data,          --          .data
			src23_channel       => cmd_xbar_demux_001_src23_channel,       --          .channel
			src23_startofpacket => cmd_xbar_demux_001_src23_startofpacket, --          .startofpacket
			src23_endofpacket   => cmd_xbar_demux_001_src23_endofpacket,   --          .endofpacket
			src24_ready         => cmd_xbar_demux_001_src24_ready,         --     src24.ready
			src24_valid         => cmd_xbar_demux_001_src24_valid,         --          .valid
			src24_data          => cmd_xbar_demux_001_src24_data,          --          .data
			src24_channel       => cmd_xbar_demux_001_src24_channel,       --          .channel
			src24_startofpacket => cmd_xbar_demux_001_src24_startofpacket, --          .startofpacket
			src24_endofpacket   => cmd_xbar_demux_001_src24_endofpacket,   --          .endofpacket
			src25_ready         => cmd_xbar_demux_001_src25_ready,         --     src25.ready
			src25_valid         => cmd_xbar_demux_001_src25_valid,         --          .valid
			src25_data          => cmd_xbar_demux_001_src25_data,          --          .data
			src25_channel       => cmd_xbar_demux_001_src25_channel,       --          .channel
			src25_startofpacket => cmd_xbar_demux_001_src25_startofpacket, --          .startofpacket
			src25_endofpacket   => cmd_xbar_demux_001_src25_endofpacket,   --          .endofpacket
			src26_ready         => cmd_xbar_demux_001_src26_ready,         --     src26.ready
			src26_valid         => cmd_xbar_demux_001_src26_valid,         --          .valid
			src26_data          => cmd_xbar_demux_001_src26_data,          --          .data
			src26_channel       => cmd_xbar_demux_001_src26_channel,       --          .channel
			src26_startofpacket => cmd_xbar_demux_001_src26_startofpacket, --          .startofpacket
			src26_endofpacket   => cmd_xbar_demux_001_src26_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component system_0_cmd_xbar_mux
		port map (
			clk                 => clk_50,                                --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component system_0_cmd_xbar_mux
		port map (
			clk                 => clk_50,                                --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_002 : component system_0_cmd_xbar_mux
		port map (
			clk                 => clk_50,                                --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_002_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_002_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_002_src_data,             --          .data
			src_channel         => cmd_xbar_mux_002_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_002_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_002_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src2_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src2_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src2_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src2_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src2_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src2_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src2_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src2_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src2_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src2_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src2_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src2_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_003 : component system_0_cmd_xbar_mux
		port map (
			clk                 => clk_50,                                --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_003_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_003_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_003_src_data,             --          .data
			src_channel         => cmd_xbar_mux_003_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_003_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_003_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src3_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src3_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src3_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src3_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src3_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src3_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src3_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src3_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src3_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src3_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src3_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src3_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_004 : component system_0_cmd_xbar_mux
		port map (
			clk                 => clk_50,                                --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => cmd_xbar_mux_004_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_004_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_004_src_data,             --          .data
			src_channel         => cmd_xbar_mux_004_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_004_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_004_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src4_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src4_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src4_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src4_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src4_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src4_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src4_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src4_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src4_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src4_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src4_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src4_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component system_0_rsp_xbar_demux
		port map (
			clk                => clk_50,                             --       clk.clk
			reset              => rst_controller_001_reset_out_reset, -- clk_reset.reset
			sink_ready         => id_router_src_ready,                --      sink.ready
			sink_channel       => id_router_src_channel,              --          .channel
			sink_data          => id_router_src_data,                 --          .data
			sink_startofpacket => id_router_src_startofpacket,        --          .startofpacket
			sink_endofpacket   => id_router_src_endofpacket,          --          .endofpacket
			sink_valid(0)      => id_router_src_valid,                --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,          --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,          --          .valid
			src0_data          => rsp_xbar_demux_src0_data,           --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,        --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket,  --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,    --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,          --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,          --          .valid
			src1_data          => rsp_xbar_demux_src1_data,           --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,        --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket,  --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket     --          .endofpacket
		);

	rsp_xbar_demux_001 : component system_0_rsp_xbar_demux
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,           --      sink.ready
			sink_channel       => width_adapter_001_src_channel,         --          .channel
			sink_data          => width_adapter_001_src_data,            --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_002 : component system_0_rsp_xbar_demux
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_002_src_ready,               --      sink.ready
			sink_channel       => id_router_002_src_channel,             --          .channel
			sink_data          => id_router_002_src_data,                --          .data
			sink_startofpacket => id_router_002_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_002_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_002_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_002_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_002_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_002_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_002_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_002_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_002_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_002_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_003 : component system_0_rsp_xbar_demux
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_003_src_ready,           --      sink.ready
			sink_channel       => width_adapter_003_src_channel,         --          .channel
			sink_data          => width_adapter_003_src_data,            --          .data
			sink_startofpacket => width_adapter_003_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_003_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_003_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_003_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_003_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_003_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_003_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_003_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_003_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_003_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_004 : component system_0_rsp_xbar_demux
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_004_src_ready,               --      sink.ready
			sink_channel       => id_router_004_src_channel,             --          .channel
			sink_data          => id_router_004_src_data,                --          .data
			sink_startofpacket => id_router_004_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_004_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_004_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_004_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_004_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_004_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_004_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_004_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_004_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_004_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_004_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_005 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_005_src_ready,               --      sink.ready
			sink_channel       => id_router_005_src_channel,             --          .channel
			sink_data          => id_router_005_src_data,                --          .data
			sink_startofpacket => id_router_005_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_005_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_005_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_005_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_005_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_005_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_005_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_005_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_006 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_006_src_ready,               --      sink.ready
			sink_channel       => id_router_006_src_channel,             --          .channel
			sink_data          => id_router_006_src_data,                --          .data
			sink_startofpacket => id_router_006_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_006_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_006_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_006_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_006_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_006_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_006_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_006_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_007 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_007_src_ready,               --      sink.ready
			sink_channel       => id_router_007_src_channel,             --          .channel
			sink_data          => id_router_007_src_data,                --          .data
			sink_startofpacket => id_router_007_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_007_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_007_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_007_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_007_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_007_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_007_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_007_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_008 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_008_src_ready,               --      sink.ready
			sink_channel       => id_router_008_src_channel,             --          .channel
			sink_data          => id_router_008_src_data,                --          .data
			sink_startofpacket => id_router_008_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_008_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_008_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_008_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_008_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_008_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_008_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_008_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_009 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_009_src_ready,               --      sink.ready
			sink_channel       => id_router_009_src_channel,             --          .channel
			sink_data          => id_router_009_src_data,                --          .data
			sink_startofpacket => id_router_009_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_009_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_009_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_009_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_009_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_009_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_009_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_009_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_010 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_010_src_ready,               --      sink.ready
			sink_channel       => id_router_010_src_channel,             --          .channel
			sink_data          => id_router_010_src_data,                --          .data
			sink_startofpacket => id_router_010_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_010_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_010_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_010_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_010_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_010_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_011 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_011_src_ready,               --      sink.ready
			sink_channel       => id_router_011_src_channel,             --          .channel
			sink_data          => id_router_011_src_data,                --          .data
			sink_startofpacket => id_router_011_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_011_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_011_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_011_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_011_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_011_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_012 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_012_src_ready,               --      sink.ready
			sink_channel       => id_router_012_src_channel,             --          .channel
			sink_data          => id_router_012_src_data,                --          .data
			sink_startofpacket => id_router_012_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_012_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_012_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_012_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_012_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_012_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_013 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_013_src_ready,               --      sink.ready
			sink_channel       => id_router_013_src_channel,             --          .channel
			sink_data          => id_router_013_src_data,                --          .data
			sink_startofpacket => id_router_013_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_013_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_013_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_013_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_013_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_013_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_014 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_014_src_ready,               --      sink.ready
			sink_channel       => id_router_014_src_channel,             --          .channel
			sink_data          => id_router_014_src_data,                --          .data
			sink_startofpacket => id_router_014_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_014_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_014_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_014_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_014_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_014_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_015 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_015_src_ready,               --      sink.ready
			sink_channel       => id_router_015_src_channel,             --          .channel
			sink_data          => id_router_015_src_data,                --          .data
			sink_startofpacket => id_router_015_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_015_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_015_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_015_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_015_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_015_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_016 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_016_src_ready,               --      sink.ready
			sink_channel       => id_router_016_src_channel,             --          .channel
			sink_data          => id_router_016_src_data,                --          .data
			sink_startofpacket => id_router_016_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_016_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_016_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_016_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_016_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_016_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_017 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_017_src_ready,               --      sink.ready
			sink_channel       => id_router_017_src_channel,             --          .channel
			sink_data          => id_router_017_src_data,                --          .data
			sink_startofpacket => id_router_017_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_017_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_017_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_017_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_017_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_017_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_018 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_018_src_ready,               --      sink.ready
			sink_channel       => id_router_018_src_channel,             --          .channel
			sink_data          => id_router_018_src_data,                --          .data
			sink_startofpacket => id_router_018_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_018_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_018_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_018_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_018_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_018_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_018_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_018_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_018_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_019 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_019_src_ready,               --      sink.ready
			sink_channel       => id_router_019_src_channel,             --          .channel
			sink_data          => id_router_019_src_data,                --          .data
			sink_startofpacket => id_router_019_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_019_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_019_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_019_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_019_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_019_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_019_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_019_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_019_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_020 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_020_src_ready,               --      sink.ready
			sink_channel       => id_router_020_src_channel,             --          .channel
			sink_data          => id_router_020_src_data,                --          .data
			sink_startofpacket => id_router_020_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_020_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_020_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_020_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_020_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_020_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_020_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_020_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_020_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_021 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_021_src_ready,               --      sink.ready
			sink_channel       => id_router_021_src_channel,             --          .channel
			sink_data          => id_router_021_src_data,                --          .data
			sink_startofpacket => id_router_021_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_021_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_021_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_021_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_021_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_021_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_021_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_021_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_021_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_022 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_022_src_ready,               --      sink.ready
			sink_channel       => id_router_022_src_channel,             --          .channel
			sink_data          => id_router_022_src_data,                --          .data
			sink_startofpacket => id_router_022_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_022_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_022_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_022_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_022_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_022_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_022_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_022_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_022_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_023 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => width_adapter_005_src_ready,           --      sink.ready
			sink_channel       => width_adapter_005_src_channel,         --          .channel
			sink_data          => width_adapter_005_src_data,            --          .data
			sink_startofpacket => width_adapter_005_src_startofpacket,   --          .startofpacket
			sink_endofpacket   => width_adapter_005_src_endofpacket,     --          .endofpacket
			sink_valid(0)      => width_adapter_005_src_valid,           --          .valid
			src0_ready         => rsp_xbar_demux_023_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_023_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_023_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_023_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_023_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_023_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_024 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_024_src_ready,               --      sink.ready
			sink_channel       => id_router_024_src_channel,             --          .channel
			sink_data          => id_router_024_src_data,                --          .data
			sink_startofpacket => id_router_024_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_024_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_024_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_024_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_024_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_024_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_024_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_024_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_024_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_025 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_025_src_ready,               --      sink.ready
			sink_channel       => id_router_025_src_channel,             --          .channel
			sink_data          => id_router_025_src_data,                --          .data
			sink_startofpacket => id_router_025_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_025_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_025_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_025_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_025_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_025_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_025_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_025_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_025_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux_026 : component system_0_rsp_xbar_demux_005
		port map (
			clk                => clk_50,                                --       clk.clk
			reset              => rst_controller_002_reset_out_reset,    -- clk_reset.reset
			sink_ready         => id_router_026_src_ready,               --      sink.ready
			sink_channel       => id_router_026_src_channel,             --          .channel
			sink_data          => id_router_026_src_data,                --          .data
			sink_startofpacket => id_router_026_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_026_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_026_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_026_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_026_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_026_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_026_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_026_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_026_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component system_0_rsp_xbar_mux
		port map (
			clk                 => clk_50,                                --       clk.clk
			reset               => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			sink2_ready         => rsp_xbar_demux_002_src0_ready,         --     sink2.ready
			sink2_valid         => rsp_xbar_demux_002_src0_valid,         --          .valid
			sink2_channel       => rsp_xbar_demux_002_src0_channel,       --          .channel
			sink2_data          => rsp_xbar_demux_002_src0_data,          --          .data
			sink2_startofpacket => rsp_xbar_demux_002_src0_startofpacket, --          .startofpacket
			sink2_endofpacket   => rsp_xbar_demux_002_src0_endofpacket,   --          .endofpacket
			sink3_ready         => rsp_xbar_demux_003_src0_ready,         --     sink3.ready
			sink3_valid         => rsp_xbar_demux_003_src0_valid,         --          .valid
			sink3_channel       => rsp_xbar_demux_003_src0_channel,       --          .channel
			sink3_data          => rsp_xbar_demux_003_src0_data,          --          .data
			sink3_startofpacket => rsp_xbar_demux_003_src0_startofpacket, --          .startofpacket
			sink3_endofpacket   => rsp_xbar_demux_003_src0_endofpacket,   --          .endofpacket
			sink4_ready         => rsp_xbar_demux_004_src0_ready,         --     sink4.ready
			sink4_valid         => rsp_xbar_demux_004_src0_valid,         --          .valid
			sink4_channel       => rsp_xbar_demux_004_src0_channel,       --          .channel
			sink4_data          => rsp_xbar_demux_004_src0_data,          --          .data
			sink4_startofpacket => rsp_xbar_demux_004_src0_startofpacket, --          .startofpacket
			sink4_endofpacket   => rsp_xbar_demux_004_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component system_0_rsp_xbar_mux_001
		port map (
			clk                  => clk_50,                                --       clk.clk
			reset                => rst_controller_001_reset_out_reset,    -- clk_reset.reset
			src_ready            => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid            => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data             => rsp_xbar_mux_001_src_data,             --          .data
			src_channel          => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket    => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket      => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready          => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid          => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel        => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data           => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket  => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket    => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready          => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid          => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel        => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data           => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket  => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket    => rsp_xbar_demux_001_src1_endofpacket,   --          .endofpacket
			sink2_ready          => rsp_xbar_demux_002_src1_ready,         --     sink2.ready
			sink2_valid          => rsp_xbar_demux_002_src1_valid,         --          .valid
			sink2_channel        => rsp_xbar_demux_002_src1_channel,       --          .channel
			sink2_data           => rsp_xbar_demux_002_src1_data,          --          .data
			sink2_startofpacket  => rsp_xbar_demux_002_src1_startofpacket, --          .startofpacket
			sink2_endofpacket    => rsp_xbar_demux_002_src1_endofpacket,   --          .endofpacket
			sink3_ready          => rsp_xbar_demux_003_src1_ready,         --     sink3.ready
			sink3_valid          => rsp_xbar_demux_003_src1_valid,         --          .valid
			sink3_channel        => rsp_xbar_demux_003_src1_channel,       --          .channel
			sink3_data           => rsp_xbar_demux_003_src1_data,          --          .data
			sink3_startofpacket  => rsp_xbar_demux_003_src1_startofpacket, --          .startofpacket
			sink3_endofpacket    => rsp_xbar_demux_003_src1_endofpacket,   --          .endofpacket
			sink4_ready          => rsp_xbar_demux_004_src1_ready,         --     sink4.ready
			sink4_valid          => rsp_xbar_demux_004_src1_valid,         --          .valid
			sink4_channel        => rsp_xbar_demux_004_src1_channel,       --          .channel
			sink4_data           => rsp_xbar_demux_004_src1_data,          --          .data
			sink4_startofpacket  => rsp_xbar_demux_004_src1_startofpacket, --          .startofpacket
			sink4_endofpacket    => rsp_xbar_demux_004_src1_endofpacket,   --          .endofpacket
			sink5_ready          => rsp_xbar_demux_005_src0_ready,         --     sink5.ready
			sink5_valid          => rsp_xbar_demux_005_src0_valid,         --          .valid
			sink5_channel        => rsp_xbar_demux_005_src0_channel,       --          .channel
			sink5_data           => rsp_xbar_demux_005_src0_data,          --          .data
			sink5_startofpacket  => rsp_xbar_demux_005_src0_startofpacket, --          .startofpacket
			sink5_endofpacket    => rsp_xbar_demux_005_src0_endofpacket,   --          .endofpacket
			sink6_ready          => rsp_xbar_demux_006_src0_ready,         --     sink6.ready
			sink6_valid          => rsp_xbar_demux_006_src0_valid,         --          .valid
			sink6_channel        => rsp_xbar_demux_006_src0_channel,       --          .channel
			sink6_data           => rsp_xbar_demux_006_src0_data,          --          .data
			sink6_startofpacket  => rsp_xbar_demux_006_src0_startofpacket, --          .startofpacket
			sink6_endofpacket    => rsp_xbar_demux_006_src0_endofpacket,   --          .endofpacket
			sink7_ready          => rsp_xbar_demux_007_src0_ready,         --     sink7.ready
			sink7_valid          => rsp_xbar_demux_007_src0_valid,         --          .valid
			sink7_channel        => rsp_xbar_demux_007_src0_channel,       --          .channel
			sink7_data           => rsp_xbar_demux_007_src0_data,          --          .data
			sink7_startofpacket  => rsp_xbar_demux_007_src0_startofpacket, --          .startofpacket
			sink7_endofpacket    => rsp_xbar_demux_007_src0_endofpacket,   --          .endofpacket
			sink8_ready          => rsp_xbar_demux_008_src0_ready,         --     sink8.ready
			sink8_valid          => rsp_xbar_demux_008_src0_valid,         --          .valid
			sink8_channel        => rsp_xbar_demux_008_src0_channel,       --          .channel
			sink8_data           => rsp_xbar_demux_008_src0_data,          --          .data
			sink8_startofpacket  => rsp_xbar_demux_008_src0_startofpacket, --          .startofpacket
			sink8_endofpacket    => rsp_xbar_demux_008_src0_endofpacket,   --          .endofpacket
			sink9_ready          => rsp_xbar_demux_009_src0_ready,         --     sink9.ready
			sink9_valid          => rsp_xbar_demux_009_src0_valid,         --          .valid
			sink9_channel        => rsp_xbar_demux_009_src0_channel,       --          .channel
			sink9_data           => rsp_xbar_demux_009_src0_data,          --          .data
			sink9_startofpacket  => rsp_xbar_demux_009_src0_startofpacket, --          .startofpacket
			sink9_endofpacket    => rsp_xbar_demux_009_src0_endofpacket,   --          .endofpacket
			sink10_ready         => rsp_xbar_demux_010_src0_ready,         --    sink10.ready
			sink10_valid         => rsp_xbar_demux_010_src0_valid,         --          .valid
			sink10_channel       => rsp_xbar_demux_010_src0_channel,       --          .channel
			sink10_data          => rsp_xbar_demux_010_src0_data,          --          .data
			sink10_startofpacket => rsp_xbar_demux_010_src0_startofpacket, --          .startofpacket
			sink10_endofpacket   => rsp_xbar_demux_010_src0_endofpacket,   --          .endofpacket
			sink11_ready         => rsp_xbar_demux_011_src0_ready,         --    sink11.ready
			sink11_valid         => rsp_xbar_demux_011_src0_valid,         --          .valid
			sink11_channel       => rsp_xbar_demux_011_src0_channel,       --          .channel
			sink11_data          => rsp_xbar_demux_011_src0_data,          --          .data
			sink11_startofpacket => rsp_xbar_demux_011_src0_startofpacket, --          .startofpacket
			sink11_endofpacket   => rsp_xbar_demux_011_src0_endofpacket,   --          .endofpacket
			sink12_ready         => rsp_xbar_demux_012_src0_ready,         --    sink12.ready
			sink12_valid         => rsp_xbar_demux_012_src0_valid,         --          .valid
			sink12_channel       => rsp_xbar_demux_012_src0_channel,       --          .channel
			sink12_data          => rsp_xbar_demux_012_src0_data,          --          .data
			sink12_startofpacket => rsp_xbar_demux_012_src0_startofpacket, --          .startofpacket
			sink12_endofpacket   => rsp_xbar_demux_012_src0_endofpacket,   --          .endofpacket
			sink13_ready         => rsp_xbar_demux_013_src0_ready,         --    sink13.ready
			sink13_valid         => rsp_xbar_demux_013_src0_valid,         --          .valid
			sink13_channel       => rsp_xbar_demux_013_src0_channel,       --          .channel
			sink13_data          => rsp_xbar_demux_013_src0_data,          --          .data
			sink13_startofpacket => rsp_xbar_demux_013_src0_startofpacket, --          .startofpacket
			sink13_endofpacket   => rsp_xbar_demux_013_src0_endofpacket,   --          .endofpacket
			sink14_ready         => rsp_xbar_demux_014_src0_ready,         --    sink14.ready
			sink14_valid         => rsp_xbar_demux_014_src0_valid,         --          .valid
			sink14_channel       => rsp_xbar_demux_014_src0_channel,       --          .channel
			sink14_data          => rsp_xbar_demux_014_src0_data,          --          .data
			sink14_startofpacket => rsp_xbar_demux_014_src0_startofpacket, --          .startofpacket
			sink14_endofpacket   => rsp_xbar_demux_014_src0_endofpacket,   --          .endofpacket
			sink15_ready         => rsp_xbar_demux_015_src0_ready,         --    sink15.ready
			sink15_valid         => rsp_xbar_demux_015_src0_valid,         --          .valid
			sink15_channel       => rsp_xbar_demux_015_src0_channel,       --          .channel
			sink15_data          => rsp_xbar_demux_015_src0_data,          --          .data
			sink15_startofpacket => rsp_xbar_demux_015_src0_startofpacket, --          .startofpacket
			sink15_endofpacket   => rsp_xbar_demux_015_src0_endofpacket,   --          .endofpacket
			sink16_ready         => rsp_xbar_demux_016_src0_ready,         --    sink16.ready
			sink16_valid         => rsp_xbar_demux_016_src0_valid,         --          .valid
			sink16_channel       => rsp_xbar_demux_016_src0_channel,       --          .channel
			sink16_data          => rsp_xbar_demux_016_src0_data,          --          .data
			sink16_startofpacket => rsp_xbar_demux_016_src0_startofpacket, --          .startofpacket
			sink16_endofpacket   => rsp_xbar_demux_016_src0_endofpacket,   --          .endofpacket
			sink17_ready         => rsp_xbar_demux_017_src0_ready,         --    sink17.ready
			sink17_valid         => rsp_xbar_demux_017_src0_valid,         --          .valid
			sink17_channel       => rsp_xbar_demux_017_src0_channel,       --          .channel
			sink17_data          => rsp_xbar_demux_017_src0_data,          --          .data
			sink17_startofpacket => rsp_xbar_demux_017_src0_startofpacket, --          .startofpacket
			sink17_endofpacket   => rsp_xbar_demux_017_src0_endofpacket,   --          .endofpacket
			sink18_ready         => rsp_xbar_demux_018_src0_ready,         --    sink18.ready
			sink18_valid         => rsp_xbar_demux_018_src0_valid,         --          .valid
			sink18_channel       => rsp_xbar_demux_018_src0_channel,       --          .channel
			sink18_data          => rsp_xbar_demux_018_src0_data,          --          .data
			sink18_startofpacket => rsp_xbar_demux_018_src0_startofpacket, --          .startofpacket
			sink18_endofpacket   => rsp_xbar_demux_018_src0_endofpacket,   --          .endofpacket
			sink19_ready         => rsp_xbar_demux_019_src0_ready,         --    sink19.ready
			sink19_valid         => rsp_xbar_demux_019_src0_valid,         --          .valid
			sink19_channel       => rsp_xbar_demux_019_src0_channel,       --          .channel
			sink19_data          => rsp_xbar_demux_019_src0_data,          --          .data
			sink19_startofpacket => rsp_xbar_demux_019_src0_startofpacket, --          .startofpacket
			sink19_endofpacket   => rsp_xbar_demux_019_src0_endofpacket,   --          .endofpacket
			sink20_ready         => rsp_xbar_demux_020_src0_ready,         --    sink20.ready
			sink20_valid         => rsp_xbar_demux_020_src0_valid,         --          .valid
			sink20_channel       => rsp_xbar_demux_020_src0_channel,       --          .channel
			sink20_data          => rsp_xbar_demux_020_src0_data,          --          .data
			sink20_startofpacket => rsp_xbar_demux_020_src0_startofpacket, --          .startofpacket
			sink20_endofpacket   => rsp_xbar_demux_020_src0_endofpacket,   --          .endofpacket
			sink21_ready         => rsp_xbar_demux_021_src0_ready,         --    sink21.ready
			sink21_valid         => rsp_xbar_demux_021_src0_valid,         --          .valid
			sink21_channel       => rsp_xbar_demux_021_src0_channel,       --          .channel
			sink21_data          => rsp_xbar_demux_021_src0_data,          --          .data
			sink21_startofpacket => rsp_xbar_demux_021_src0_startofpacket, --          .startofpacket
			sink21_endofpacket   => rsp_xbar_demux_021_src0_endofpacket,   --          .endofpacket
			sink22_ready         => rsp_xbar_demux_022_src0_ready,         --    sink22.ready
			sink22_valid         => rsp_xbar_demux_022_src0_valid,         --          .valid
			sink22_channel       => rsp_xbar_demux_022_src0_channel,       --          .channel
			sink22_data          => rsp_xbar_demux_022_src0_data,          --          .data
			sink22_startofpacket => rsp_xbar_demux_022_src0_startofpacket, --          .startofpacket
			sink22_endofpacket   => rsp_xbar_demux_022_src0_endofpacket,   --          .endofpacket
			sink23_ready         => rsp_xbar_demux_023_src0_ready,         --    sink23.ready
			sink23_valid         => rsp_xbar_demux_023_src0_valid,         --          .valid
			sink23_channel       => rsp_xbar_demux_023_src0_channel,       --          .channel
			sink23_data          => rsp_xbar_demux_023_src0_data,          --          .data
			sink23_startofpacket => rsp_xbar_demux_023_src0_startofpacket, --          .startofpacket
			sink23_endofpacket   => rsp_xbar_demux_023_src0_endofpacket,   --          .endofpacket
			sink24_ready         => rsp_xbar_demux_024_src0_ready,         --    sink24.ready
			sink24_valid         => rsp_xbar_demux_024_src0_valid,         --          .valid
			sink24_channel       => rsp_xbar_demux_024_src0_channel,       --          .channel
			sink24_data          => rsp_xbar_demux_024_src0_data,          --          .data
			sink24_startofpacket => rsp_xbar_demux_024_src0_startofpacket, --          .startofpacket
			sink24_endofpacket   => rsp_xbar_demux_024_src0_endofpacket,   --          .endofpacket
			sink25_ready         => rsp_xbar_demux_025_src0_ready,         --    sink25.ready
			sink25_valid         => rsp_xbar_demux_025_src0_valid,         --          .valid
			sink25_channel       => rsp_xbar_demux_025_src0_channel,       --          .channel
			sink25_data          => rsp_xbar_demux_025_src0_data,          --          .data
			sink25_startofpacket => rsp_xbar_demux_025_src0_startofpacket, --          .startofpacket
			sink25_endofpacket   => rsp_xbar_demux_025_src0_endofpacket,   --          .endofpacket
			sink26_ready         => rsp_xbar_demux_026_src0_ready,         --    sink26.ready
			sink26_valid         => rsp_xbar_demux_026_src0_valid,         --          .valid
			sink26_channel       => rsp_xbar_demux_026_src0_channel,       --          .channel
			sink26_data          => rsp_xbar_demux_026_src0_data,          --          .data
			sink26_startofpacket => rsp_xbar_demux_026_src0_startofpacket, --          .startofpacket
			sink26_endofpacket   => rsp_xbar_demux_026_src0_endofpacket    --          .endofpacket
		);

	width_adapter : component system_0_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 101,
			IN_PKT_RESPONSE_STATUS_L      => 100,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 102,
			OUT_PKT_ADDR_H                => 42,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 51,
			OUT_PKT_BYTE_CNT_L            => 49,
			OUT_PKT_TRANS_COMPRESSED_READ => 43,
			OUT_PKT_BURST_SIZE_H          => 57,
			OUT_PKT_BURST_SIZE_L          => 55,
			OUT_PKT_RESPONSE_STATUS_H     => 83,
			OUT_PKT_RESPONSE_STATUS_L     => 82,
			OUT_PKT_TRANS_EXCLUSIVE       => 48,
			OUT_PKT_BURST_TYPE_H          => 59,
			OUT_PKT_BURST_TYPE_L          => 58,
			OUT_ST_DATA_W                 => 84,
			ST_CHANNEL_W                  => 27,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_50,                             --       clk.clk
			reset                => rst_controller_001_reset_out_reset, -- clk_reset.reset
			in_valid             => cmd_xbar_mux_001_src_valid,         --      sink.valid
			in_channel           => cmd_xbar_mux_001_src_channel,       --          .channel
			in_startofpacket     => cmd_xbar_mux_001_src_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_001_src_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_mux_001_src_ready,         --          .ready
			in_data              => cmd_xbar_mux_001_src_data,          --          .data
			out_endofpacket      => width_adapter_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_src_data,             --          .data
			out_channel          => width_adapter_src_channel,          --          .channel
			out_valid            => width_adapter_src_valid,            --          .valid
			out_ready            => width_adapter_src_ready,            --          .ready
			out_startofpacket    => width_adapter_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                               -- (terminated)
		);

	width_adapter_001 : component system_0_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 42,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 51,
			IN_PKT_BYTE_CNT_L             => 49,
			IN_PKT_TRANS_COMPRESSED_READ  => 43,
			IN_PKT_BURSTWRAP_H            => 54,
			IN_PKT_BURSTWRAP_L            => 52,
			IN_PKT_BURST_SIZE_H           => 57,
			IN_PKT_BURST_SIZE_L           => 55,
			IN_PKT_RESPONSE_STATUS_H      => 83,
			IN_PKT_RESPONSE_STATUS_L      => 82,
			IN_PKT_TRANS_EXCLUSIVE        => 48,
			IN_PKT_BURST_TYPE_H           => 59,
			IN_PKT_BURST_TYPE_L           => 58,
			IN_ST_DATA_W                  => 84,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 101,
			OUT_PKT_RESPONSE_STATUS_L     => 100,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 102,
			ST_CHANNEL_W                  => 27,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_50,                              --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_001_src_valid,             --      sink.valid
			in_channel           => id_router_001_src_channel,           --          .channel
			in_startofpacket     => id_router_001_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_001_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_001_src_ready,             --          .ready
			in_data              => id_router_001_src_data,              --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_002 : component system_0_width_adapter_002
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 101,
			IN_PKT_RESPONSE_STATUS_L      => 100,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 102,
			OUT_PKT_ADDR_H                => 33,
			OUT_PKT_ADDR_L                => 9,
			OUT_PKT_DATA_H                => 7,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 8,
			OUT_PKT_BYTEEN_L              => 8,
			OUT_PKT_BYTE_CNT_H            => 42,
			OUT_PKT_BYTE_CNT_L            => 40,
			OUT_PKT_TRANS_COMPRESSED_READ => 34,
			OUT_PKT_BURST_SIZE_H          => 48,
			OUT_PKT_BURST_SIZE_L          => 46,
			OUT_PKT_RESPONSE_STATUS_H     => 74,
			OUT_PKT_RESPONSE_STATUS_L     => 73,
			OUT_PKT_TRANS_EXCLUSIVE       => 39,
			OUT_PKT_BURST_TYPE_H          => 50,
			OUT_PKT_BURST_TYPE_L          => 49,
			OUT_ST_DATA_W                 => 75,
			ST_CHANNEL_W                  => 27,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_50,                              --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_mux_003_src_valid,          --      sink.valid
			in_channel           => cmd_xbar_mux_003_src_channel,        --          .channel
			in_startofpacket     => cmd_xbar_mux_003_src_startofpacket,  --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_003_src_endofpacket,    --          .endofpacket
			in_ready             => cmd_xbar_mux_003_src_ready,          --          .ready
			in_data              => cmd_xbar_mux_003_src_data,           --          .data
			out_endofpacket      => width_adapter_002_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_002_src_data,          --          .data
			out_channel          => width_adapter_002_src_channel,       --          .channel
			out_valid            => width_adapter_002_src_valid,         --          .valid
			out_ready            => width_adapter_002_src_ready,         --          .ready
			out_startofpacket    => width_adapter_002_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_003 : component system_0_width_adapter_003
		generic map (
			IN_PKT_ADDR_H                 => 33,
			IN_PKT_ADDR_L                 => 9,
			IN_PKT_DATA_H                 => 7,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 8,
			IN_PKT_BYTEEN_L               => 8,
			IN_PKT_BYTE_CNT_H             => 42,
			IN_PKT_BYTE_CNT_L             => 40,
			IN_PKT_TRANS_COMPRESSED_READ  => 34,
			IN_PKT_BURSTWRAP_H            => 45,
			IN_PKT_BURSTWRAP_L            => 43,
			IN_PKT_BURST_SIZE_H           => 48,
			IN_PKT_BURST_SIZE_L           => 46,
			IN_PKT_RESPONSE_STATUS_H      => 74,
			IN_PKT_RESPONSE_STATUS_L      => 73,
			IN_PKT_TRANS_EXCLUSIVE        => 39,
			IN_PKT_BURST_TYPE_H           => 50,
			IN_PKT_BURST_TYPE_L           => 49,
			IN_ST_DATA_W                  => 75,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 101,
			OUT_PKT_RESPONSE_STATUS_L     => 100,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 102,
			ST_CHANNEL_W                  => 27,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_50,                              --       clk.clk
			reset                => rst_controller_001_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_003_src_valid,             --      sink.valid
			in_channel           => id_router_003_src_channel,           --          .channel
			in_startofpacket     => id_router_003_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_003_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_003_src_ready,             --          .ready
			in_data              => id_router_003_src_data,              --          .data
			out_endofpacket      => width_adapter_003_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_003_src_data,          --          .data
			out_channel          => width_adapter_003_src_channel,       --          .channel
			out_valid            => width_adapter_003_src_valid,         --          .valid
			out_ready            => width_adapter_003_src_ready,         --          .ready
			out_startofpacket    => width_adapter_003_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	width_adapter_004 : component system_0_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 60,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 69,
			IN_PKT_BYTE_CNT_L             => 67,
			IN_PKT_TRANS_COMPRESSED_READ  => 61,
			IN_PKT_BURSTWRAP_H            => 72,
			IN_PKT_BURSTWRAP_L            => 70,
			IN_PKT_BURST_SIZE_H           => 75,
			IN_PKT_BURST_SIZE_L           => 73,
			IN_PKT_RESPONSE_STATUS_H      => 101,
			IN_PKT_RESPONSE_STATUS_L      => 100,
			IN_PKT_TRANS_EXCLUSIVE        => 66,
			IN_PKT_BURST_TYPE_H           => 77,
			IN_PKT_BURST_TYPE_L           => 76,
			IN_ST_DATA_W                  => 102,
			OUT_PKT_ADDR_H                => 42,
			OUT_PKT_ADDR_L                => 18,
			OUT_PKT_DATA_H                => 15,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 17,
			OUT_PKT_BYTEEN_L              => 16,
			OUT_PKT_BYTE_CNT_H            => 51,
			OUT_PKT_BYTE_CNT_L            => 49,
			OUT_PKT_TRANS_COMPRESSED_READ => 43,
			OUT_PKT_BURST_SIZE_H          => 57,
			OUT_PKT_BURST_SIZE_L          => 55,
			OUT_PKT_RESPONSE_STATUS_H     => 83,
			OUT_PKT_RESPONSE_STATUS_L     => 82,
			OUT_PKT_TRANS_EXCLUSIVE       => 48,
			OUT_PKT_BURST_TYPE_H          => 59,
			OUT_PKT_BURST_TYPE_L          => 58,
			OUT_ST_DATA_W                 => 84,
			ST_CHANNEL_W                  => 27,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_50,                                 --       clk.clk
			reset                => rst_controller_002_reset_out_reset,     -- clk_reset.reset
			in_valid             => cmd_xbar_demux_001_src23_valid,         --      sink.valid
			in_channel           => cmd_xbar_demux_001_src23_channel,       --          .channel
			in_startofpacket     => cmd_xbar_demux_001_src23_startofpacket, --          .startofpacket
			in_endofpacket       => cmd_xbar_demux_001_src23_endofpacket,   --          .endofpacket
			in_ready             => cmd_xbar_demux_001_src23_ready,         --          .ready
			in_data              => cmd_xbar_demux_001_src23_data,          --          .data
			out_endofpacket      => width_adapter_004_src_endofpacket,      --       src.endofpacket
			out_data             => width_adapter_004_src_data,             --          .data
			out_channel          => width_adapter_004_src_channel,          --          .channel
			out_valid            => width_adapter_004_src_valid,            --          .valid
			out_ready            => width_adapter_004_src_ready,            --          .ready
			out_startofpacket    => width_adapter_004_src_startofpacket,    --          .startofpacket
			in_command_size_data => "000"                                   -- (terminated)
		);

	width_adapter_005 : component system_0_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 42,
			IN_PKT_ADDR_L                 => 18,
			IN_PKT_DATA_H                 => 15,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 17,
			IN_PKT_BYTEEN_L               => 16,
			IN_PKT_BYTE_CNT_H             => 51,
			IN_PKT_BYTE_CNT_L             => 49,
			IN_PKT_TRANS_COMPRESSED_READ  => 43,
			IN_PKT_BURSTWRAP_H            => 54,
			IN_PKT_BURSTWRAP_L            => 52,
			IN_PKT_BURST_SIZE_H           => 57,
			IN_PKT_BURST_SIZE_L           => 55,
			IN_PKT_RESPONSE_STATUS_H      => 83,
			IN_PKT_RESPONSE_STATUS_L      => 82,
			IN_PKT_TRANS_EXCLUSIVE        => 48,
			IN_PKT_BURST_TYPE_H           => 59,
			IN_PKT_BURST_TYPE_L           => 58,
			IN_ST_DATA_W                  => 84,
			OUT_PKT_ADDR_H                => 60,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 69,
			OUT_PKT_BYTE_CNT_L            => 67,
			OUT_PKT_TRANS_COMPRESSED_READ => 61,
			OUT_PKT_BURST_SIZE_H          => 75,
			OUT_PKT_BURST_SIZE_L          => 73,
			OUT_PKT_RESPONSE_STATUS_H     => 101,
			OUT_PKT_RESPONSE_STATUS_L     => 100,
			OUT_PKT_TRANS_EXCLUSIVE       => 66,
			OUT_PKT_BURST_TYPE_H          => 77,
			OUT_PKT_BURST_TYPE_L          => 76,
			OUT_ST_DATA_W                 => 102,
			ST_CHANNEL_W                  => 27,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_50,                              --       clk.clk
			reset                => rst_controller_002_reset_out_reset,  -- clk_reset.reset
			in_valid             => id_router_023_src_valid,             --      sink.valid
			in_channel           => id_router_023_src_channel,           --          .channel
			in_startofpacket     => id_router_023_src_startofpacket,     --          .startofpacket
			in_endofpacket       => id_router_023_src_endofpacket,       --          .endofpacket
			in_ready             => id_router_023_src_ready,             --          .ready
			in_data              => id_router_023_src_data,              --          .data
			out_endofpacket      => width_adapter_005_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_005_src_data,          --          .data
			out_channel          => width_adapter_005_src_channel,       --          .channel
			out_valid            => width_adapter_005_src_valid,         --          .valid
			out_ready            => width_adapter_005_src_ready,         --          .ready
			out_startofpacket    => width_adapter_005_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component system_0_irq_mapper
		port map (
			clk           => clk_50,                             --       clk.clk
			reset         => rst_controller_001_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,           -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,           -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,           -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,           -- receiver3.irq
			receiver4_irq => irq_mapper_receiver4_irq,           -- receiver4.irq
			receiver5_irq => irq_mapper_receiver5_irq,           -- receiver5.irq
			receiver6_irq => irq_mapper_receiver6_inv,           -- receiver6.irq
			receiver7_irq => irq_mapper_receiver7_inv,           -- receiver7.irq
			receiver8_irq => irq_mapper_receiver8_irq,           -- receiver8.irq
			sender_irq    => cpu_0_d_irq_irq                     --    sender.irq
		);

	reset_n_ports_inv <= not reset_n;

	sdram_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_write;

	sdram_0_s1_translator_avalon_anti_slave_0_read_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_read;

	sdram_0_s1_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sdram_0_s1_translator_avalon_anti_slave_0_byteenable;

	epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write_ports_inv <= not epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_write;

	epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read_ports_inv <= not epcs_controller_epcs_control_port_translator_avalon_anti_slave_0_read;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_write;

	jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read_ports_inv <= not jtag_uart_0_avalon_jtag_slave_translator_avalon_anti_slave_0_read;

	uart_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not uart_0_s1_translator_avalon_anti_slave_0_write;

	uart_0_s1_translator_avalon_anti_slave_0_read_ports_inv <= not uart_0_s1_translator_avalon_anti_slave_0_read;

	timer_0_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_0_s1_translator_avalon_anti_slave_0_write;

	timer_1_s1_translator_avalon_anti_slave_0_write_ports_inv <= not timer_1_s1_translator_avalon_anti_slave_0_write;

	led_red_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_red_s1_translator_avalon_anti_slave_0_write;

	led_green_s1_translator_avalon_anti_slave_0_write_ports_inv <= not led_green_s1_translator_avalon_anti_slave_0_write;

	button_pio_s1_translator_avalon_anti_slave_0_write_ports_inv <= not button_pio_s1_translator_avalon_anti_slave_0_write;

	sd_dat_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sd_dat_s1_translator_avalon_anti_slave_0_write;

	sd_cmd_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sd_cmd_s1_translator_avalon_anti_slave_0_write;

	sd_clk_s1_translator_avalon_anti_slave_0_write_ports_inv <= not sd_clk_s1_translator_avalon_anti_slave_0_write;

	isp1362_hc_translator_avalon_anti_slave_0_chipselect_ports_inv <= not isp1362_hc_translator_avalon_anti_slave_0_chipselect;

	isp1362_hc_translator_avalon_anti_slave_0_write_ports_inv <= not isp1362_hc_translator_avalon_anti_slave_0_write;

	isp1362_hc_translator_avalon_anti_slave_0_read_ports_inv <= not isp1362_hc_translator_avalon_anti_slave_0_read;

	isp1362_dc_translator_avalon_anti_slave_0_chipselect_ports_inv <= not isp1362_dc_translator_avalon_anti_slave_0_chipselect;

	isp1362_dc_translator_avalon_anti_slave_0_write_ports_inv <= not isp1362_dc_translator_avalon_anti_slave_0_write;

	isp1362_dc_translator_avalon_anti_slave_0_read_ports_inv <= not isp1362_dc_translator_avalon_anti_slave_0_read;

	dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv <= not dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;

	dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv <= not dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_write;

	dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv <= not dm9000a_avalon_slave_0_translator_avalon_anti_slave_0_read;

	sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect_ports_inv <= not sram_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;

	sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write_ports_inv <= not sram_0_avalon_slave_0_translator_avalon_anti_slave_0_write;

	sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read_ports_inv <= not sram_0_avalon_slave_0_translator_avalon_anti_slave_0_read;

	sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable_ports_inv <= not sram_0_avalon_slave_0_translator_avalon_anti_slave_0_byteenable;

	motor_cw_s1_translator_avalon_anti_slave_0_write_ports_inv <= not motor_cw_s1_translator_avalon_anti_slave_0_write;

	motor_ccw_s1_translator_avalon_anti_slave_0_write_ports_inv <= not motor_ccw_s1_translator_avalon_anti_slave_0_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_002_reset_out_reset_ports_inv <= not rst_controller_002_reset_out_reset;

	irq_mapper_receiver6_inv <= not isp1362_hc_irq_irq;

	irq_mapper_receiver7_inv <= not isp1362_dc_irq_irq;

end architecture rtl; -- of system_0
