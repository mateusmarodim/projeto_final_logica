// Copyright (C) 1991-2013 Altera Corporation
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs for
// use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
// ALTERA_TIMESTAMP:Thu Jun 13 12:38:48 PDT 2013
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ihUGOGOz02u4lqbSQOMupE2NPYTnrpmIFIqN9zBDqM3SbYZB6hxx2wZJ8Z0eo3LX
0pzCaySonkHq8PL+NFwBBKkfU9LXJDEJMMMAxpt965NRwIg3oLpJYDwblCHFlTAT
441nxK9aDX9zwRk+2cQdjlL+iohXSwBR9rJ0Gp2wO8Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17312)
CMaeveWz/NhqFMJaCID3DLUIwWrxGVw1Y1FrEnErVT8vNbjTvgTyGjsIfHRgGMZx
twjL0xYokZJt9oNVsbK9fmnrVwVgBmKYjOlE+JObtWa+JnCGvGjtcuyfsf/XTIgo
7wUUJu69M2PsN/ZrKQKQm3sPW2ijRV/bABN67jo2Ba4KpLVNJzxxPVxS87SBW3m0
e9LTlHDdUE95HME5w4aaZm94aUKyn3gD/mw/eGYoZqfR+Ds08QeqL2DtSvPnkJkb
lWIXdszRo/nlGvYI60KAn/LEXPmTciE0nzGrlAv8zf6CpSfxILW+AeIUYXRdfV6/
xOjD+a6mnuSI0B/501/imIf0MRzYpsj6KZOwjHigs0bzpAkcIIqfN16vFmxU6qPK
emeRTBCXqwmOAHgln7SG7Vu33OD36O89Z/9lziyCHB+eXxDUfWJ8rfEHUKy0W5gd
xSJi3mZE8WxfyX8fSlhjnWLFH2lQAejxPX9BFKuHshk68NPCf7sUyXY3oa0MR3F/
0JDdRE7DC79/9rTAv4mFXwEncOrNP/amdBwcJYdQtVRgjc9Y/TrylqOUytUuXvZZ
agUrKsf5A3ueF0rMDUNGG0vKqs2JVYC0PFiLeWK8k02nldslYhWIDb6gBCZUomWb
OFnJjZbBdvuHRQo1BUvkP54I6PpqCeIcjDxIWt7Oy4ED+Cau3nUYu7ALkeZVDLb7
9kd/QjMrtLfKKpS+ogB+tw74wkuGIXymeL468k+t6oSumnlnjRFOM67zRFnM/QoN
So4AX9HQVU0BH7NmLpq3EYG56q6fSVtpZpgySDexE2lratiwZvZLpL+RoYJfFD74
Felk9IaovHMcJViEnOksbm81GcChedG6YT6waRsxZs7M79X/B1PDAYYwh3s4q3XJ
MMSfoV0MNp+dCmWwnVBx86NfJlFfnNchKg6PoXTP/9RYhrQPDop7+3rK7W+Y0+7X
eK9hOXOrXmyQJifew7HxU+kMiaBsHcl/WqlAIcYfVx9eM2cUlawlFAahABSqNPml
jBxNS2zXXf5gem3o87GcA2/cP9sYRZtWDr/s0LOI00Z9o6qVSk1k7Oxaoi0oZQiB
7S/FBJ5xxu4B+sStbmfN8mSxL7Lqh3WLbp/QsK9g2O5fhUpqybcfqd0VpgjHmIfs
jC5gBR3D+QpDyaQE1yankoTawRYSbh2n16d3uUx6W3oEsx1MuPzOtMy3BsZoeP/1
kSHZKFTpWxKnhkVYhpqT2gLuoLMj3FYyGF+5jJcjYnOEwB7gj82gBCcUPBKekXur
75HC1Hmi5JmUEC/j7RKJpCdw77lkKWUlNljo68CvixI1aSmK1u2PhArapkT4g6Vd
j4ljRhToYu6uDh7YrBDFSoB6q7t3Uhlq085axaHaLaUDhNmoy7ii0XpDrJEC0Iv7
5UXF12v6RY/Xh0Qt7fyhyCKeqv7rzh3SftbgU/36EHhv5ht6veKFU4ezTxo6Zt/0
E57nGIqTyLG4vDmBu7lpQVKGBh7vwwKeWMuEOD4MCxdZNhY/30dZ7Sbzw0KvdV8L
/1NkORSuMjGbJl4xMWLYcRvdOEIVLtSi+srMWxftQ8ulPNW0gsvNJPd9zZWZk1HW
JnHGstqXwfjHcJaGwvDBl4h+a1FXFaDXGn0d7pZSIzpdLJtJZdjTj2RRzDxmSNHk
irVRLGkl7H2TI1kQudVHO5n5L0WDSEhjubLmZcQ9C5bQndVt4NUq6CWvgbFP4jCt
+XHngHYqtLi31B2EOGtO7oJ8NZ62XP8Jq5ESMECo7eSGX+hl6j9Nsrf5a/P++vcs
0roBsy1iJ7+KBO8zN0GKomDH1cRWOrzhquBJs2NZF2+/jJXjK+/WwXpqpP7o9U6w
Q5V4Myd0xvIcOQx+1t5Mt7ezc4HncUxxakaLNHRP+neNCajLIgmk9UL7AJOqCQCJ
GTacGdcsnUAu6rDayj6JQoCdbIyxkFl2HPlQx9nnPFOQA+IxzC5+iFqBjHsNywOz
cKfkiap4bdrr29dy+ATZfDDvxn37q0PEfwXL7ZGhbs00pL7vCUeyAdPuj2fQYkqx
LbqKwvM4MAh+b/dFggObLerjnb0h6IBWnJUfdomkJKOa3mQjlV+BBoZxgWmKAIVm
2NzkZ4302WLcFtBEtOguZNnysFoAgOWRsYiAT5Z4uDEVf3dQDUHMViNYNhufP41O
HojTt2FEmq66Rqw4+U1Tun7zYlNOHM4zZWHTrDcrD/d3teduVymb2Ka9AqvkzCh9
rvwmNRixZ9shOfF/HdbkIZFDsEiJX3hZO7ZZrNHKWIzaxbCGTVO28ZDcXb9hSaku
4+HEHrNpBYiMg/nLqXG3Ln48IxHkYRJthkq2/aS46A5Im0AU84BvZN7W01hY/TzD
AQdxQn5Ja1/8Ksg5B8I1AUP/KtuXaParY5LXbYVIVTKFGoAS8kkzwM7gG/ual4Ly
TFpd0DUPHJXWn9LOuFlk+tbisPVYFWC08grDc1Ur06YwVykpqC7yLFAF3jHF5D5q
Trgk07x/x7Bc86v8O76GbRlvR2ZqxLNz8bRFYn2BkOppTM0KdS9fMABORjZ8v3U5
kw2cApA6HUDGcVGxsH9JM6yZeJC3qZjQtG8Ug61kV5i+mJ3KqCYazWwNbhnejpG9
gk7nBcc00IP85xOmiy1Mm3otGD7I6nGB0ULXW1oBfifCuQdgceRKWfKDlHJ8dgdS
DCt/Tw13/YzbpuoDqbHiQ/qOdBEHg0vmG2ywvVG/idhdn267TclOhmAkSIoXn9g5
QxjdE/Ox9Q5aIk4aZz9nrProe8IhaJgbyLbjdkjaFwHy6ROIHOuKcyr0dGdqYUCd
5TRIezZGjf4eO19+UJlmabIs0CMdeqz4pT1gMIknZKQZ7nRbea/cBJ6hsHxfAaHj
Sg4rkmvcKdSux0ssyAliaM1eRL1Hdn8W0AkEEeEfacgA00beA39F9O101u2S5j5k
/ZqtOo49s2ofuD5tEwYNdbqOTvqxUCx66xcJ7QlRp7bjEFBfNTs9nmTLoczulPVe
dm9I9PrbaHn0Gl3RnGVUbDO0dBX3/3leu7D69AxVsPyxrKpASy7+hOt9BQPouxiQ
CLUr6V8pF4i072wcYBMJuNN2smoGFiJY3cjCqju4uDn32JZZX4lIdmomUNuF1LLD
WZJrdgrprEMJ4khFb4dB8ccdN8zbF4evGIOyb3gBYwXP4RcdCsEXOx08UV2bNLLV
Vypv6s7aFSacW+ISZeFLW9jyUgTPe8QyXumsnk4X0brnTPH4uturK6V5Dx0zYOn0
lsyB+vdLrqI4UWwKJuoT+E8oKw6BSUVubAP+FWSdiIh2ZxlrVrBCxIW4YAR8IRVa
DcdslgfF8tr4uweWCZlqMF5oMBb8DClZcG60sZJpwhLnZd8EyDzvfqLVcPN4QaW3
FHgHD+lwrZ4vWGpe1clLuE2forpEtlIVwBYvH2vrY1/nOwBeE2nMVGtKWtBU5D/K
aqBSlOEHWwqWa5TrSaIq0+RZdXuYmngXthxSjFr67+oKkj5cn+I0pZ/eaXRe9zhs
fFMGxzKwgJadN1uK9gcrdbPWekOeIOnsCASLQzga/ADaAmPKtQLFGX2CwBKTODW6
P23HDNeZ0drHjAP2E0xtAs2/mp713/APL6lj/N6P+YoHT82/++TdownmCQUqkY+N
4R0+bsHqiap02PiCz6hP722H+OkFTuTIl67+2Z6xTzcRN5RK1z6nhJ17zzVA+ool
dkyLJ561llHB0Pp0O1VxXM27yTw2cg/tMFXicV3qwsN0Y4ezSsPnt4kU+s+cAs99
0qCMOlRtTfUmzyfUHc9acfmKbm0+inEKZHPSuMiE3U9Ys/L0KMifif3bMzOo4dSc
HLngB3rY2YJ+AecwuoUd48LK1Pxm8b4WHzc8dddTXhsoOiYaIIKZcWxO6wOL/e72
SVyVr8dd2JA4zs/J6I2HXCI+TQyll1y4R/vGLpkvFAlfRasSGH5+5y3uuQoAOQFI
OFv51M4KTJ2Er5n7wLOLdcJUd6MGJeZrHvxIT0eo+lixmjZg4lJ8f9I/rdbTP73H
qMJh/L2Cn1MWdJTt5Ih0EyI99/HXrk3rMitILAyupCtS3lqf5/HhgI4/AYuN708d
KRYWOQdQjkRGu5P+2ghcmC6l79UINSaBHRCbOmUGHQzBd/xM3NyhkdUDMGJ51jaU
R7XQSftlTpc5yWrn2QoswHaQEecc6LvQ76ef0uWVx8S63B3jQGMDwmK/X3Vgk4O1
NzXRsnjw4qviPwAMXQ0U4gQ14cT6B6nlzIkKT9vsxMdfje+UUI+gHzeqhfThgXRO
2E6glF6HOXM2kG8oMqnS7fYiL5ZT01hCXYWrtXxsMEfUmQtGiQe5ahrGd0SmnNSS
EIQlzUsarz3U7iotYLJPNjsINbRQnc65WXLLIlWDxtlKIis9225Spv5MNSF8m6eN
FBoh7U9uYjLe6i1IAWMx++s3pfsb6IKy38UF+MU8SyVIcnlmamlslEAWHZc0I8ol
01TRuVKQrQZ7elHX/hnoMFTtPtad7G34Kwq4wvtMNA0xfXOtB2Ta3hy3FD1eV1jS
vSK7DSkTQyrkPkuezvzEZCRh7PUZMcij/6lQTTeb8S9XJDzKfNh/Z1v4/dg1juE0
P3ZjvAcLPX2fZMfFb2Mc4mKUYKMeA0dH0A+pSGJGQ5NqeC+obOhEdH0SgLU/MGZr
Cy2VcVjuVBxi38D+BeqzsNKLM7jAgH+dcJymIwMtopnrKKPY1JkmGKWe9SM5iftm
7UZE8yGOH4FZjbLPJRoeM1LX0nivPSWTr8Qz68g07RE0LdKtgr5b+vH3fu+xWxeS
JwnT6yneDx6020teVBP+9YJFQhRgS/eeQaJwX7afc31xu+3oxyh2vFWuAjpv8Jpj
/Uo+2vsnn7FJD8EOLmmOT/ZxYoZv5QyQ1PLzNy7QJRqczlOTb/jg9g2ImAJkqEwM
9O++AMbcmoadXm7AH2HvFvUUCJ4FJ05HUQXn48+9gqqTH/iYyCCsJ2yCKmjxpRFH
nLmBjRaDGOM30uPqcSa377OGxktBKpMD5uH992CgcinGRl2k/S5nRBo7piurQdZy
BxJkzeoqj+hBdfankxSOMC5fZ2383HY8x5vh/v1sCqOyD7g9jazPOnoyQib2bjI/
GHZ/rehptj1jAOjk3IaPLC/UkNfnhNZ86XkXtGVrA1sNVnSEJk+NtQTavCuCLGQu
H0mIcweB/2y9jD4whb3rsvG1WTsPzL0ThR43gCRgVHq3+3YN8EUeM59AMEKlZX8f
70Ds/YdEYWL+CBO3SezhaPBIyAUJkNFItBbQeyVXy29ekllwyQCjScU2VW8EC/xr
+EmyUKqU5Xe0DzicnXLscfOQv4M3PurvjaW7MyfaKHPkqqJwgYOAEq987FaP56pF
/N8hPCltc0nWhZXbooRTgAXakUjwSo7WmP921HHpnTVSqm6I/Rv5Ua2kMCOvwq20
JqJjn7AGkMS8ftk00X7ea3S+09zkX51WuNtgRmUcF/1lKAlUdeY7Ydudgg83k5H6
AImV/cXq7TRENbT4ndbSw7AdqS+BranQDeiOSljhgrkDdvxuxqEIDBk8AUYWTBqK
UQN74sBApfF8kFNYE+IqW/Wg6IYQawApd/1aTMcxzv6WpcfDfb8Qy8BddnyTGMBT
cDE476sqo/vgH7sjwNOJSPCsnINghA8lcDAwRN4Nb9t5VlSS2TNoJctGinFWWVQm
DUgbIUQldNkx1W8H+1UxUJclBx6UB1H1Ml2Th9BNByubKxPcLaEIGKRh7l8MYxwf
KElPgx47REt0xS/BM4+GeVM4pCY199fj6dHhs8qohj8lmN5FTDz3xGY5xbvg/jdR
WwawAGKSJwKMymp+gukoLQTyjN9a15qkMs30AU5fCsw2b7Izdcebr88pd7lQ4Lph
MMdLTdddS8cG+x4mLkM6giFx+amt4djJcTu5nHWxf1gqAc5jgK3pxZEHUW67GVCC
NVb1SMSRHtbQlD0hXjezq0lAk+G0r3J6O9pEk6AWyT2MpVDn8GBFplZV8mibNojY
HdYB8pQCt2cSNyWfdqsXHa/Y0Pyu42jiHl6vJ7hkIPD+JJhNp6ojCUfEvNzFczCj
v+V+vT/P0F+qs9XNhkg9Uh1T2DWPPMCrmI/Ua8fOE+VdIY/Ex9lrYWI8vt0EglgZ
De+1o9F1Lzkh5Hh/81QUQmtIAO06Jg21hSPS62EWHciTCouWZm08T5WHsBSzi5br
g2Ua1FLIptmTZyAFUG8WvIOjHyxk2Orry6KUbarMq4DO2knvEDbcHicZ5Lk4zmJ/
0i8685s9iQdwhRa3jgxAKeTDC+TB0ZGAT75MqooW6ba8SqUjUHzxOlwWiTYAY8kf
pRdF3M7KU/9aawFRQoVG4/KwmMKRkRGwbciHl9ZgEBfLzvrk6vVKqtCLemgfrSNb
kxAWO5efvM5lCipEnTr6YvwjpPExlz6crQG6K8Lx0/gPNzQXA88IoctjBf+1Yl7r
bkcBii8Y/2RsitSOm8eeuLRRhEs7E3oolVjITWpTuto8G8tqAuNPaOhbnQTCufBQ
vTmUUmRUzVepsbVG4oq4dzch/5KzAYrhndrSXvRpaboiZKbH2Y7W4A0rkYcOC8vZ
GRsQdw68VOQx29kW9rBgGU8zUxH1ftsAQ0heJeRn20jDlekD01MPcT8zqDmLdR0H
5GD2nqePNcU776GLIrPL6H/YRQOIGWzyGESOiTPABbHjA3huXPJe8yYYjcSVpWxM
ycIXGBTZykqDT/DmjQct0x0p2MnHzx2n+DLn45wNIJQCP0agf2gWI5e9iNbDK4S0
CpX8sD6wYNRH/VbNw7Y6ypoCgN9uZwGhY5gSDG2cDsiq6Q52AoytXPmc7I3Abbzz
+cDRvFp3Iy3JhqaPUTnwaPKSRuajGyyj1JHoqgRXjU2Oa5fw9CUSQDYbBwmc7/6N
ASqOpemKk4TwRw9W6ogxFiTp45o3SyXFBBkmDbrSHntFutRyUL9OAPF9mVIOT07L
xMgJ8ib3NVUHsuDaG4XtSlCE1hZUacZfBn+y+d85iz5/XyFFupV1fNoHZr7kyI8/
GAQOvPxtTmWAUHQjRVTWQowzvqwVZxTdT4xf+OFWEeCxg2mGtUdyh7ysH5ZN0QQi
WAlh7In7gvVTJpxAfFpPGUjoJfDgpSQl79figlcIGsDb9uNnAmlh2Hhvbm9UBYlc
JJNkhfbSkyw0iUJTWn8H6sb32KEFH29mWJS+U1/9+ovaAtK6Gr+wAodAVICbhcXU
/SvDA3LvyL+MgSKLlQ2N8rPxayw4ycSe4W742MVgD4v32b7CjFolhvcTcbPGidMc
5jpzaHPpcxeYe2PZJXxt0OFy2GyHN35sPwesYMrmCUwZhtaPanFkEvNOjkCG5zBz
19zN6XYaLnDV1ma7Gunwp08I9kmHY1U/otgc284Wg/IejDI+16rp2UxTMQ04RCd7
Yk648pcTU6TI3gv3uFCd0euABEYCpNNr096NxYjudsHHHZecEuASDbpJTvxnlUmW
DUPCsOd5F94xcRuBK8+IYRIx/oCS3Zyjv3vnBeoq6icNIIGBsUILsgv0we75FJNL
whrYViuD8g8EXYtWBIIdIyV5BQkDQvE9NNs6ImiL60feCPjTnmqYwGNRKRaOmoqt
kVLQuGKwvlKJAenFxy1t9yhRnj0d+6PcCu/KBfZb4CA6TIFRtgRVj98IArkZuSMd
WkmPNelkQdE9dRZI9vc6pmJHtQeiif4N50UchFo97JvTDEKXzSYO96aSPIRJRehm
uUQsufMsWSs4aqHb6rGxmue3OEAD2GRhL6JqhvwWP0HdMhuCkg7Q0rRFKiabc8cP
W+46Dhfi76Lo9+lp1kmVfodOdoyFZd6+nsFaOBirbLwspMxZKbzeZYuPmWE+y2iD
5mW6KFL3FbFfLQRTUAXheSHS0RJefvvjaDWDVr9Vk1fmOdj3WOLPRTpx9LuvybCl
iIX9SJM9UMprGLa2poayVQg381Ys3/p3Oqxj/u4VhWR8av1gMpwhvjvlhzEke7fj
0D+iaOPoY9waJjpt6V0dNPrlwJ78XFZ+SW6TEPiLVULcPK9osoLAdq84G/TR5Gby
Tl5DaxX1ySkwx0DAquDBiUAfizT+H6jF0KnlDOR1+hYRR6N0XDzSX/10ytV1TEOg
GPO/MMkFfyh6xo2OqTJnnf8SInW4BiS4uCbyGW2luHlWolifq1a6U9IKFCaoK7w2
l+MiCLuGkRRm0gHf6S20EogbdbQc+kFm7E15wBMzTIuuHEpe6v1TSZVYma03wcwK
LOr8HWfbXNHIJtyadQFJCK29uabjbWWgROpECTaRLj0jH40BUj2VDOW42ZHfU1Yn
+tX6fyOEZBWD0So1QW4hnIEYeZLUxLeJupxmtaJtOm/6mwNrzAVCkjJcMk9dS0U1
Q1vKv9oMZbZh2TzM+bm61q3suZVv8PG9imzEQ3RfLnE0y3MHuwwU0DBvkbr9gnRd
mudlUUv7JBdgUC4mzHYg7FURvt+J+YLOcZwyukh1Aa1++7rSTtHWAjmpP5OAkLvn
/WSiA0UMGtwbphxH/IRtOkkPO4wQ5zkMvOHmacHym0ywBqUIDI6RONnzyaKRsU/q
997GVhRpRQTcowQGgbwRmezcIbCQ91zWMU5jWVOBhU9Sx59RwcIaMiXTES/kYnck
2nZ1vQ72AW4yiwRV/vFUr2Uh8qfkPj8P7QcpYleU0Z4IyDlkNLpU7oypVyPzHzhb
w3xX4EXsfcKoqh7JIYtAawVzlm0ng+NO6hDL/fzYjtFdCUYDHtbiWlvCtu+n4hY0
HiZ0Kr2yrfxzKKp01xR7WPxqt8gunredVNcyWH+iwHqIM5z7aOBDLQw05tErEVYX
W81IDU6Jm0HAT4Hjf2f698IqGcIzmTnolkTJhhpPDGE9fixGOBxGALEqbxJE3gw/
QYPIgLC3xkC1p4at7zTVFdK7fB/nASjNjTDkM/TMJqV2Xsk97OhkuIHZRs5WN2Vj
hWBaZUfsV/vnvSNGNd/9kotRLVDWu184LBJvx6XD2p7+n8IZyWidNTiCEhrKN7Q2
QrWaoNVdJ4OuylDbF2p/oJ94t5mHfl+ggTEGlDmWE9SNJzAVY8cdmTH+0hKQF+/g
zpVne9OlEUhCqP0xc6pc0XnGaIYN/RJLRgfvCKhXYRQD+DCDgJLNXIeVP3CjWWzz
3f9P7xNprSuSvjWIDfwEe/pYBDpz1tDjmtC7ZpHyO3UQov72qWI3rx3lpdk+wtd9
w4HSymJA8P4SBkuJI2ZAlX34W7gJc7sgM5hMfQ0vmIcltwqtgNL3cXGHigEOeS47
xbhtcYxF3+yBNYi6hFxKcCqL+le9tjxlFza/1loTjSLCgV3JkdYjPsN6MAM0mdTJ
OY2Pf8rr3KotZcb7Nvt/vHh4TJ3GrmDRtBM66xpmRpfCqLdCp6IK7zf9mRQgiDKc
z3df09e3QjFeZq0MbAJxRxQZxO690StMq3KV3poIt192qnU+K8JBTggEeOEbDjRq
kM04+1joERh9TstmBLUxVfFirWHg/bObVjwcZqtqSQCOH1/SoDCUhPqAcOZ2n8oT
pEo1AHy3XGmUERpadZmnUvJi0/E6H03CSH1XitXs6ww2u5/szagNIUM52wad49oc
cAP7RvVzCohBVEAAAn0WffwF/MQcIfyWsanoUhMzazQShNJZK4Lco9CLGWgOKBRS
CS5WYC7BMVt8TfvH5GaQs8zRTB8zIdBm5/DQ9S9xDVCVPSq2pFiovvl848y+RGQN
QqbWEJSmuHDhOrDLpr3VuYLSeib6iao91o8kGJr60VCpGKmlMaHoc6n0jPadYyYh
8DTN9rnSrltsOwniAT6v6dq5768uE7DSoyfFycAnSwfbDLN/CiP0K4k3jxGHk+gK
0N0L5I5rEvyL2OxjXx+TIxFY+CchEMBOs29QXx0fqDikZkzkmuYVBvyUC/bsJxUz
rzT8+lZfQSGAwHSJFLutbcSegk/DI/n99CsDJb/s+vgj5DK9+LJBhdBtLmlPLkgm
8yQRBDwh94+lBliHxtZHPZIIJBbTHa5j+RwuSK5zW6aRKoNbae48u69T1OItr9LH
RCWC/IQSshTVqBVmujvWREbfFhwMfQZVSwi2MUrI5OIsCObCWoYzHizPC03UHg3X
pt2t/77dsurUDtfpXronMq57CnPw9B9fSOLItDdQmedHwdyODknBdA2dtEODFSbd
AtvmTsNJG9DLtzIA9h1yfUjz9V5buNMxCcRTn+dUVYTY00x30w0fs7SM+ZDgb4VV
LeDV/DU1qY36lokXcqOpZly95BfnNvPJAmV8EJYsGNi/EPuTKFgvxaZU7VewuV1h
MlD3K/mqPODmO4mAeSBM96HSL7Klm2D9CKIGhMpQLvV7w2zhgfBoSRxPQxX98tah
TUQPxhO+wg7zBhZ9mgnhZKl2ptdTbZTpzZZNRucO4uj1BDAlqazv+9orAp8jdotx
OPEcO1t4lxZA0y5ymxSAt9ra+CdP6jKWfyNyosA/DenBNjZyI+WYUKMfcYz3Kp41
1ix6lEqahSr3YSUzQPH7eWkvIhCkQpHDFkw6DjrGlVmpsANHNFfkHMqITiAQQR+N
VOYawySjVTHkjxZEU1nfO+K+zPSp6Mk7gCzihEtALGGZnQSHdK9d3JNGqLidxN3W
ULi5PTNH8gidrjLwXnPOgNMT/eYl/6LSVHtt1wc/lcugm4cyEGHbbO+VXUUAT2dn
Kmt0X+/09fTQAtwf4zBVGcSEaYnd56DksZH4w9igFCLPjrB53PXQWI2gN+a8/3r8
ryykWsOO7hctlqvFk7uDt6W72V330i6XBgLm7ptrdAFrzqi5LKnPG8Oq/xcIJwn0
FZ3Z2QBrNExV38Z28numbJdR4HGmB2GmxxXgrPluN/W3siDIM9p/OWD4USWRYVet
YGWDPLj40QJItMlpzHDjzs0f8MNfDxDTwLb3LFbmnlYHO31colUGuXvGXKUMAyVX
8fU9vPw16cW0u6cRsx3pguJI+D/6D4Ms01RIHCb/0NmWgKr6I6qtiUrLIiMnsIvV
BruIPlMKz7r4K3iF15VHIDdnx7JUwkZhFASwLXuo/QMikDFcXM+qhKdnP8RPul9i
bliDxUKYSivSjY5Wg7MBirFqZA5xjRlmnIK/IZNzSUWAFX+ENu89aEn8xNEwCP5n
UuPZ/QtvujI5XYJt4VwFHM49Yif4MUw01JFadMmU27FgIloJAPeq/yz+Pv0oLqCc
gQHpuvRtrYRKGuJZHVWQcRwcGaZl6Cw70rZLIuZcFswB+BWSDJqLk3ldRXuLChtr
GQPJWsJDbS5I0PaIf3JuhIk09MjGzVl9PVUMowQ1r1NrAkntBrqEny3C+0LNhaXj
GpseCllsUaykOAW3X0M8jKRmaNQvdCDZiacjIKFtSX+mdkUtiy9vAu/reSMPgSYM
KTpTWm/HvB++Sq0zmSVgckCVHshPKSXrG0UflaQr7xuS5+EGuY5jQk2K/m+cHzGa
jpfv/GLLuMybKdCdKYydIiyUfnz5nOaI2XdPb8YLEStpL7WtZ6fZNIMIO6zTgOtA
e2hJBFltBFjJtGxmBf6kGfVbVxLEN/WtNaPrnNBcNDTg9MpYLnq+PSUT8kH2PFbv
1IOyXzIvOQyEuX1EWc3SjEL/MvnoJxCiKPtCIMQLy0AwCPRerkKokKaoceziQ6YR
mA71wrmDovuK+W+Tz3hBelr1Yl2XgCMN3RA5fW7zJHWYxpfN8nrds0vdG0H7+zcU
6c5PoH+ySARO0X8eH1v0YuBGH0cfJ1ryt0eUhHw04zcs7oJHxc4beiCiaEtTUoaL
L5Mse+jaZAXKvjZZpzXL28OKxGKfGC1P5+EsMOWEk4AcfTMX5VlkiLgFDP9X0N68
R0RtAOr96U+iAKPdwXrqSxsO+1skkQidSj0Er74e0O2LRTXrM486J3xwS7ICCNNN
yD+n/e6PL5SFQwLi35yJv10BV3b/0ZJaf1Ydo0WJ6rqJr/gU84JCkvGMFAunbCAv
IUp0RG42ixk1CZde7aUj41J9LQuqV0JaTq4qnglCStEA+/1pbNfwqNtTEvVFSGeb
JmwN0WR+D0dueFoQu4d8JDfIY73wZlEGqN6YRR4ANI+K9IwaIiIIRRSpG+pMxCM1
n3A3yXKQ7cdifCizXYUf8fVY06fV2s+NAC09B6YI6hD7hVLWgh2chWk6mkfVQEXg
tLyof0b2ecINKsEC0pQ+rsnHZBkjlwxMD2l8ixuMwjA7zN8koVZJ7NQu0dNBIpP2
EKKSDiGFFKawsV3ZIByoPLawkeccw7QlX6fwLFaKfl+c8i2N7X/8DHjPHCoBdrL7
DTIhbflwM+ZUjYjClTnMROAnfEGd1b6ATlnBVdGPt7U/vLJuErvnEFgHqKRv0qjb
6tH9MFh7X4afdUVmoCAJ1CYCBbxC9CtilopZ2vFufWBGdYtl3uiBSt3bArcRZdfK
jRg+LqEjSZxhU24uOQV19JUvJGFHAxJjj+MRlDPHkle+n2fsNxVwaIH1ZmZZLrUg
ct+W7H9vP87D+vyL1xOwjBffpNj16ZxXYnIz5vDrzhUfGhZZFlWnAJ5KvbQHPu51
skEkREYE5a8TboxsReLgATbFh/FitxuYeb7NIAzXH+v2HfDA+4t0zDMdpDcQV/uQ
9pG0nJnCd3Qn3VyrvIyIdOgHKZDfRmgyTlvkBUKZqwLzmmxK98s8DZkBHc5useP8
Y+1Of8OLXMRpMNbXKNA8+7WTF0qAxjYUeJY1iY2fUjXoq/jwBSN/LiiAvm5jLiYp
xAm0Qu1KffebsI38uUk2YIRdT+lXomftz+SGpgQMLr6rmqAQml21kjhxQrvALlYp
v+hdhYnmYKOYlCyWZuVMPfPJJRAKPVJdQj9vUQmwKIlnHalLB5JRKIcCVIU77ABP
DmGYRYzfdYF3Wtgv60mkIBmT5tk8fiZCmq/QgtoeM1a4fnod0yPD5uarTVpFuf+B
0nIHrCYnzDpOSUGBKWB145wwo3adsMd01SNwPEgqADz5ad/oaDQLsMgLmdrookwu
V2xDERRPK5BMbJE/jC1+gM6sHkmjUQD6Q1XdC4oPX2naJWi+rDpMth5/zEzwXWo7
2WAHsBW73ehALLUtE/UQR8BxDIhjkoCdtOa/1ZX1GqhfO7SyzOkY/z4ff8BzaqfE
6j5AejSlG5YChymdGSv8nPHC0O1E3U9K9LzFxBs45O5g5hvrquIv1r4xskvuZRWB
Bfh6aaK3XugDTB0lBBsTPel8Wo0W+Ggu9O00z6Uq5+7w+QcEhFMJy0vLkGvZMAnP
F5vUXoLCLL3oUJ8hi43dDWJFVU357H+8PvdFyEpmGSUl1t4ckUU/ezW64TKmdOYI
fp7678iKiagU8yMD7Z7sZbGAne8icydirEXZbHtRA3hfESE17+CRMbSUBaJOT3nf
+B0qr87nGWRKnjfOcDfQKTUnHOUjVw0vAjYCdrYONlO7LQnT3OYu6iKTlIv1XyhL
+z7EQ46LU+RsZfWXVq1PE8yNFlnejHwariq6eHbdhzguB5HvN4RJ7ntbgeE2e3lQ
MCdx6hc2GFTfPgZ1MzRRTLdG44TLNtSVaMFS1PYWyaNLs+XYd/mkmrjCu+/uWIZK
Es9IxWUlH9IA6GjcPCaTWk0mvNcAimf171MXWg2UPUKt4kD4JQg4VCgKgtUM351T
ZbjpKBLeMJHasecTLiUc1Mx3BzdbYRTDq14FZwPyV1hNj7QZnYNeUHRzvsWp7tr7
UTWxMV2AHU4MVdQPavODhqcpUfsMwdM6JAUfyxDYbc3JqRfYfsIQjXGA5VA2ppju
l8Ii+KSiEXrrVJWn0rh4UprHMncuxkZpnQQsCMAwTGzOawlGNhRBdbsdQO1aQ8Ai
v1j3wwccVYNjFgMxMZ2Fnl5DR44NuwwllbvVLRhfDo2gfv92XXw5l0PAvGWV0Goc
MuoJLVRbyOqErmw38+Kjtb/IpDD3usxpNekSScUKD+Zf/+Vn2c3NM1f7YRwrIKpw
uVOo04W9jPed7ZQ6ZghEYcYgfAhBlfry7PwFRp1FfKo1tQxgXuQlp6hHVaKUhU4F
sW7z53qyymv2OCDxPmmvVrRG0+jrJ+H++QEjSZYSMNWQOgtXodU2Uw8aXYerB6HR
T3WgiWmrBC1X5v0Ql2aIqn5/uD9vZYSp/1K4Volqz2fIf9j34hivZwM46Ghe8plX
+yXasqp6ncmLZfxtRLtJBdm0v2ntMdlq/4tOuwzNBR3/DsCq/AC8Zb6jJZcgZsJZ
wizCCHXeJ8tS724nej7SiYj0l3MR22o6dr9+I/Z5DQFzuo3mQWTlztKHKjsprq6L
nYEbvyldOCucmo2U+LmmbN1DiNvtV+j1OJFBoaIOqcfErJ//L2NT7ZwXm2ezrkMx
Nvb3xUp+9626mVrlkDxABBtLAuSZK/khLwYNkwrxS5HVoTug0gPx2rIpLNurI8o/
oj1uA3sxUXqrmIYMydKP5kuJ1IzCq+VuwghgvoYBfD7ycGGHvz/j0qwqFVE8FMYy
XkC0yViMVkxMrkqzuV3GV4HayyLQvTB66iFisj+A/GrobjKDs2s/9BBYim2yiuag
V5N+t7rPGJfLavunJ5MLVrrWqG1iUHYwhZ4nk1p7y7Ay83AEZz1KxiejffoXh4EI
KH7Jl9lr2FtnLBaZH8TUl7zQPMzfVERgau0QAwQ5M0QU8Nws6SntMZqyFxF1S2VS
ngyRg7F55mqc8NGNlkcItbsN9uN+XgG2Ax6DnnjzM7oE7oUp4Y4cFXBvi5ZNfk1P
JdW5bBI93EQwW3My8G1Gmu50RAFJsqF7igVEUaxGF02OrpP+MxfGXCaNbbtWH7hy
0SNEoVxOlqJmRMT2k2M1hvTCzAn9kR4imPdiPq0YPQuVouFNj253xw1MjjQrcY+H
d6wdhpu8ya/i9kZ0H05JOUcvbYjiidwwRpF3fWu7cn2FXm26C6uyaVG1YO68iwtm
IqXg/w4Yd2DmUgldHY34LXuhhr3VO96twZTbBXdEfFI7e6Nvq5qm6umDm++jsKeo
PozK8yhlUnTFZDjoQUvsc9geCxsjNej6eX1vZgNA0yyM5z3SBl13I5dgnCq8fwwk
CHxmRmPpNi0usZLi0ort6eAM2dRmMctlr1V9EHurOe3R3PA6Lh7VHpO1fQmBwlPj
NwnWMoVavqbYxS+eGvq0CFk2N4DToI+SztiF5J3SpHofUrrhSviSWm/JdK7vBNaa
L7FUKqpqLxgNQrJYlnKxUPbop/hN5oMAhmabVrUxd6a5/8Jv8Wiok8LdbzlydL3t
O1HAbYoe9ENRzBzcET10v95FgKVK2KM5oZnZOtg/B1DSM62asG30OsiroAviBW0b
Zk+ivoB/6KSX7bEuyguePItR4HM/yx0smKZMykU1TeyjZIqFZeCJutkRQj/9TYcF
OJbPu4i+NPNIwHvaVgUCUciEZll/cU7M24YoJR3WOcaf9MfzCm1adaWXJSoZIWsN
B/DNcAfgbcozzRtdxIX7VcYHx6qQzYD8qODwiByD0eeVKjpO3hR0Q4wjzbbvTtFi
kiLunXQCpFuujBEE4Q2nNbnAt7tvU/zLKn2yvi4q2VZ36nYJW01NyH2dKW6LkNzk
inF9WiP9aM7GUCUD60Va1fDml9Ea99klVZVTf6+orSM00XYLcAXc+kJxWM8Ywx9j
VSFMvzT9+9PUzHxVS1Y2d4ER0+grmgB/j+2XK96jNcvn5BFKlkNGCjokHfN7HPi3
MmotjfKnnsKrBJMEZwhxjIjB6SXF6kepaOZN8VZViVlA58V4eoVX/J4BHQDHWeUd
roW+GhJFKzbgi608Ens/t1VwZoSAjkTw/xarSzeNBKOyVUizgTLn/AN0OtBRSfTV
UildSFr1xqTN0+0mDxYE2tuBJSo8gqJ5HRFvYRubtWVgfM7hYCRkywtYWCyL+Kvl
Erq2n9lLTLYh27ujnovTEgltkp2wru53rglIpJ4ElqPovlsQ3DGsSvvasq+GiCU6
risnRIhlfUCJBnyI6wPN90k7WELFct7/lLMUdGsLgULaV19woWvoNDhqohkiLey9
0MlO/4pt0hINTun+8KFjc0nHRdCmkCB47AI+y52avAwRrvZIkEw0CDJ9Di6pezND
B+Aqu1aA+uFFlujdM6xoscHMdFV4KJuV10DisWwMLscy4pf49Xb5J2EdugAdLBty
zjWZj2DF9VJhKXjxLm9BSsKBI9HqeDylAOHuB0esEUJdN3S5naqm+DwN0a+TyGqq
Oa3nJEcuyqfnuYXNepp3WErb8UisFumiBVT8NmnnWlQrmnCmqD3i8cMpXm+JPE+S
aEUAoD5fFAkzcJHlBLZBIcmtG0VLPd+kDrVKRtyhPGZWcE09gnE/ldzHfYIHOgre
GyRpLoosMoOjeI9Sax+LCtsl9PwEVN23Ra0RhKD/aqGJFfGu1Ojcc1GdLNPlOFvf
YoLEjzAujAN5X5Z1QSKGL64IivKai6F0GT7p6ozgGHp6KiaeA27C1RHhJP+4hEwY
0LcdE/pvS/qES6a+fidudoE4xejmWtj4kgSfeXf49s5cVC/Shx0niVQKMZO2Dzea
aEDnShQdrPq+OQKzhgTVIJrFOGZJAZ18LO8Svf9JPF/dmDcyQZTXLGwTnmrGCwMG
2T55wvbGHHpCgzJJKaxObfhP+5qMAAoRFj6FlFegKtU86OhUYrMcryddYG9USJu0
Cz5o8MAs2uslUOtbVk1Bu4lONrWvKOZDfL3pKeVPKWJLfN3COxhRjeVZSSe4pjQR
oU3GsxqFt5ONaZ/GLpRy7Qs5pJBn5P5Lht7kIu7M7cIxfrnVdLSOt3an8slclSim
rkIJRtfgehZMjGrPL4HhYBp15JykvzCekSNUKXBmSrptlD0wc66MNhVEn+fQD6Qw
YJK0Nw9TDOBKpj77aiyR5s9HgmiGunlpuTeCuE9lf6qnCMuFpUgQp31WUXNXmwhV
Rd/UXR8DLATPIs789OUmsnlfRiu1IwbSzNxcoRS6qAXEciFockEzvvQUkAGpKby8
/sXJQbg7eFI9Rg67Qcb8VTxOBsLpjYrk5eADcFB53WnZYibCOjnW2H3Ud2BBjY9D
7lvX070DNmoar7qGl9/HQDYvdwZXl0x7FtPq1aG9mggS+aMPqI1C4LbOAqtWXE7y
tceJZb8EdQR/mIoKJsTVa4jsdtyTlfjM3I3LBqF36kpSwjEUNZUB/mJfVcdtpltt
tZ0a30GOF4u7DELcjTeuwECUYlDsJG+vJnZBatDYAK2WsdJuV3C1mHwgfVH7AdDx
Ln/o3vCGL6XaFfv02JGnhqF79I+RhOL0s6WgPB/DD1sF3/japLrwBQky6pl+wqPE
XZ9pMhNt5iVG6UVetuDnYihi+9AkTUscV5aEniqpfggObHRO+JyQmzsXB+/lWvAU
oTsDDqK2BdnIeA1WmlPO2MB5DqXXCGbFVR2J4ilcjvSP7G0G0XH+A7guvQs2xHU1
Y4tnur59O8BGHYMzDxp6S6ST2hN/RqEm8rBKsORio5ndTqpJRClRlh0JmtUAePwl
1oMYdRzXor/WgIWW2e9wqXPAJIvTtZR549NV5m52HGnQRNSwPyfYTz5ybCLXrf+R
61Q0mBYdwToqe0x8ysqK3GmUmNJ2cB2BJtHqv7XFZzQUQD1fS/a00bPNG0btd8gY
WdYjaGmCRKmfcEhbu+/m+3lYC6YFwXuCCiIZsvMOMVgH728Qy/mpyL1CgRc/N+h5
rd8RyHX/d28vjUknhOr3FF7VWi20V2wj8+Y2W6nYE3qiqrg9BG7mv2iGf3MCDFCa
M6+g2ZszhQ2Y+GQxxvAgmR8IAT+2BxL0IMho10Hzz1XNBKC1LBswPzv/Ztv8O8aZ
3R9e7sBaMecZtLZFU1306BKCgrRlpRnmrBe6z6Z3GjDLfemiW15CoYkiQBmtpPqb
EgpaFtyZCeuzBAWyFfajCK7YfPrph0yphEUqdqnfcvfn/YOV2tAodaB152HfacLt
kFYn5WuAtRbzHfpFjjvYelkR4bGXJuU4ERYdNs5JPZoDsy9yDzS2bErbYlI13ZE5
UxkT4TaBeCcEQ/dU5sY5aUfn2jUTS6M+mzP3b/RjN8ml6WVA25wiDb753/TeePdV
QUHqgLibcQpCTaonJkYb2ymPtpGIUWC988wWIzpQSzGAJG246yk6XO2nMwUGP0Cp
0p0OYWnI42AhEtetgRar/UP86CFRQ2Dv8xk/ZRkmGYQRcQZkOlPw6pbqqVn5ZTOW
vXruPicCpFZwq6vFUIIkCQ5S3Nv6sjq2mVy9YxaH+efS+lP4NlqlEhLS9RahLYfj
wXbcuD/cqPX01uPEnKou1rW88FsmSwFHsNVktyoaO+VbA3TRNa3pLa5YjpnFf8Uq
umssyj/2UEt1QsXvnuY7EMtz6jfwXEUEfU851xp9MGDbUVg4SZ7Be9m9jXCUEQ8+
53Hs5oF+zfvGqkQWmv7wT2+lvfiAX5FZkjs6A3dGVFvxjqlDteo2zK3LiLXY9AJy
qAg3RbbCkcjytrZHQ4UWYvz4j1Gc9IqDHvS5FDnb/jtxjG4O1eokmUlIfcgIkIaD
QuPIp9PvF+8XqDD5qs5hqED5y5uU4h8vYP1NpAGfRlnQHkRXO5gFsRO1XXclAj2O
BR7IKhTlw3PgsZDinZjcZBFJ4wwc7W3NkozQmhDv//KpjK+DG12Z1MG9alyGE5BC
/IhNxo5y63YMcaEnl+TsTTQw53SzaWobWRtMd2IZMBg8JdkHy5MIZauHNggjG2Ww
odbw1z2fVhGpCy4V/acD/P8siGTURlxM0iodqvL4I6xFdXtb0lUIo0T7UHQQwAkC
SiiuOeKpAj8ZUc9jIP1795tWpaYMaMT5OvOEhUnXJXzXD0X5Q2co1gteRstxbRjx
SCxk48QOHqaX0Sc79/6qxuZ36fO90Es0dWDoR7gIwEufb1Y+skn04jpVIfQbKeN0
Q48B2Xdm91VAN0AVd4ZvpfL3U0Dx7/2YVM0Rnn/tcJRnodg0s5W16CHU2cBcid3w
eNKc3eSbcPsBB6jRKyJdK0NOJyNjQlTXb9H4ulyJc6/ib87HR9Fb/cG2/eUjWwbK
qqo6v/eGjZOnxG+pGatgS3OSV/sg/1QwhL8PjCUgAS9LqWnljwGWtydIQSpFpY9B
5ElfFJx+/PMURDYd2/hJ1/b9FxYtBcofE4SMB/hzHQi0hvbevj2m3GyDrldOO4oN
N46HLxOM7S7lOYCVwsu2C61DoOrlAETiVMbzulC9MX3YiT5+IBkraAH5+x8Plqry
KQkgqE0qo8IM48aGIsNl7F6fT1fIFMeCzvBl11C8Q0YIv1Lfi8/fQrNEvSx44Bvv
ci14sOUsD+PR7XS3f5ckBK21dsq+KthJ+kqgycZnD1CPHglamKCS8AY6RaNS2jll
81IOOUsPy4T/NQVsZ1eFsp2rG19g1vUCXQojN4s7tFvpIEtOheWW8MrD6B9i/pUC
eQMB8V6xS45ZHeE4hcB3nBVZVHuH/WK7YcCGD8flmZkqWyUzvDuxCh55VWUt2bju
+Zzf8ie0yjwbDzG38e4PCLO4Ck0ChyBKvFKE0dur6y1iEQc8th7G5DzmVYRPzzAS
N9kIaLvCDu8lS8/T7JiSRELdbiud/Ana5yNXTK1tiOomyqF6VuqK+eurtvskl/7Q
AUmorjP5XoRRWY1BXOzQ/3ZzDTbEwAx7dZLQjIdUmpfvkS7z4Xl5ikZ4tsbA4SAk
X7UNM/r8HHy+h11/2+tJh7Id977qNufeghghWxSHZ0COWcM4HB1OVxAI0dfSjBVb
Rq8PJ8kLpTS6P+0hwDajiI4+9FrExPrc1nQxFIC/YMEZi/N1jrkY/jWjAL0GIyjf
rU6r4+lQe8PbIfRLwb9I6E/okE0/eu7vDdT23JVtAaRjqIZ7ehLzQofMpgxmaw1F
fsrXH7meI2FKvuDSdGNkltPv1h0+oNFHAApu4x6ghcdn/iUEGR8flcQ8svWOTsTW
7Y2LhYMqsGzG/+g/veg+RnSG0ZsJZeFnaRtCM2sEYRr9SRsdu4dSrDuBc2LvNFkk
JJsFOSW40EKdp5ugrxcNtLPlUwnwFHP+BjLGj5azItML24YHdo2ZDsJSwb4GJYNw
YSqZXTTHlhL6yLQSbEd5ZgEuNfAkUzesJ+ydkwJvQbJvnMWFwCi1UVkdxgZeRaKw
Xj8yHleV0n6O1R87D9nSdGcSeKrzk2GlSXPvq2rncm5os+g22kgr2Dv3OQqSgBeC
M2IQ+X/u4nzHzEHEhysgF8muJ8L2a9WpmjJ4dLLoB6l4sKVCYe81Mf9YtXrZwZBI
CPYaCvi8hJU2tVVHqSuLPKvDbSlzNk0pWiczXJYj5Pf+8aFxnAcaSKHTbdhE/15s
3WUvqqi9pkRqk91BcYFRnycNqlc3TU6upXwO3g5SGwmk7EOIlqRwMQxZfqTBbHD+
I7duaSrkwuOPapaTjwOpmic0LdH6+lArk0fWipOeCZ+IqcEqfDX2RaYhziIuWohX
3c+GPgnWZmsle/7LLAjw+YW444sj7KXg1OaiHZCSsUvJjIWQtOsOjY2Ebycg0OMP
RfrP9Q4dOmD1xgjlgGGETbhLiReBCNhKbd7S5hy7basKq2rg5bcNDUR7ukMz7IOt
IVCDUgUlMdL0vSi8fiayFl0smyM0QucpSUPHO2ND/UD45Dl2ZTvCbIIafvsT9bB0
q7JleX+u2H+vFvQN+KD1IFyHoH6EUQLQj8UycZZ+zjQYn0eGhDQnp8Dn3hwVQ+A1
oXejPOUEeKUON5hczQ+A7KE97gtyhhFgVy1NueEh57+frDUVKX4kjYRi9f/N7UzU
pFkDskCCoGSNU+q8j05RIGi7UcHwYiUyDgMZcwkAPuBBSK6c8pY2PYbd7Ok5WQ1O
5inmtH1LNaXrQ7C/GApDrL8bu1vBeQCFvkGrx8XsscHZLXpINTiLePVzLSCivCge
goQcHF7G+JXbHMnA//vMcu3yp7Dl5tPxCD+69e9lnnyn+z37fxgBiXUoIgOuW74k
NfctyHIMsDQ11gBnNjGVU1a7jUpr4RQZqKylNBALPVliWQiiPDv5ZrjIY55paAlj
67ByPfw96ZDL8uUrkLIS09rQUs//AD/eoa7zWoL7UH+lVYbNpQOX2nJNBaMhc4TT
VXUbuJlyXElAYJKk4heonSZHKLK2qKV6JpIDB5MynLkVFQ4xzOrNIkE9PuS12kLs
ITXxK+hA9K+u3WjeU7cMt7Cdu6StOpl0sG49lPuH6VhEbxM4cq8wHO77Wfq68IWE
SMwwjcGlGFGVl21njDwo9TutIXwqnKdIeh2TQrET/fETDgJlOkk32X6S3AcBPEB/
bJwMAYsi0TyYLAwDRyaWvR4pdfXzpT/KptoAQ83oVe/Lq2jHWZy6yrEooML4YRmk
idtp8od6sB1liFUG1MJQHZodcwrnmq5JIn0d5ygcbUfYiWsLiHru9hGmvOtbBE3I
17NK2Uwx/I5O7GdO8kP1a3bbJMFXyknfAhWbGNk1fgcvhOh/8ahGutNj0x7gPaj1
p6x6tG1qoOh0fpdNhKGK1lyhYCsWZaJTPgYlWM8NIldt1WPMcKdKRnk4lJtXvDZO
D4jnqv2rGxkm4co63l9ckqQoWBvjj4XK2rMW6ssbsCrJtxji4miezSNQGT0QND0M
ka31dTUWFpJn/yOfY1prCHb8nUYTM1v8fmyLSKkz3Fn7E0LnjddTaVKtBMY6MYAB
979PYIlp9VRuJpZZ0HozgiYQXesJM3JbssQ3l6MhBQEzHP7ORLB1RlMo98uLoBN8
1fuZ3u1ycy9dGqrgmWRitqqBLO4HOtSRrWD96QR0IeL8+l6ruk3ziadszSME+Ex5
5QN/Hh8DCorJ8DFZeouIFfxU5MIjYSZupxTxz6BjBqdzEdTiNp6I2FGtW1G5rz7l
3aF4z23OCYwhgGOhMAtgnXFiJu5QFM6M3tb3zYkYANEw9DDiJ5o64aVtckITZWiR
aUUF+OU7zru0BINJEyEUtSmTklqGQ+XPTBz2s3SCRsQo6QDKF4LZ2QlQqMkPLndR
QsM1le00CDROnSyGT2OEZnvCnxX3Qpcl23tZe9u+qK7RYUUJbaMm2mNtTfHsD4yy
4r0pxtBV58ZaI2SK+LaDcepQiZb+cKD9SVuHDNytes2x8/3h/nrhwdJYfLcw6L+o
m6spdSNHCH6uAVDgjfFyNV/UEdQaZKxqyr7+Bb803kL03Wc62S6tscoYHkEy8xCO
ic6q+uoPAWAy2et9z/3/iAKzTpDhhicgFzJBq0Xas+OvdbDWIwYrTsu58mOc2C6S
PVejC3HVo3FytlqVe1F+7Sh5v+ksm/PnbIDZraMzyW0KcjDCvcS8cCx54L/shGZu
35pIAqSDvC+yH7ZZTO5ktBMG+Ygt7VTswYYfSkMrq9lSp80u4sQhtBt4utSUAkNM
1AW38qcOz5NGfkGdmrzcW+lnDz8MtOiqt5gC7TGveRz/yNbIzej2ewd10OEvbayE
gZBHyfNJYGJVgJwhIrkJQu+TRr8Q95fCiVLBrcVWge9FmvPGYDjd4yyhmH3EsQ6L
u3YZn2segeeeESiM8XcMT+RVvtFJyBnWUJQMqcV/0uOT5LMTVq1SPc0AaS6I7bIp
FO8tikVkiWgsnELrn+v09hFD4x67AJQdIM7rxUrHu+yva+11+dceCgPCrWKWNKtQ
5h9r+FhrTLBDuh35d0t5pybU7cJzf5PepFWdEz0krP1MtcNnZXN/6GiDZqh50Eql
yAayDWNoUwYwKNzSpXKLlJCwvz21XEoPMZvwyLWf3ZGSpaDkQLWhgLERf9mS3ORI
8plF44KuZxpNMt6+hSXfyKOygM/f1AWVQZlZoYVT7n3Mr0Al9NEu3GcB5fLqF2oM
xQ6R/4woMntWFQ5zUlpM4WRfCxtX1wSpGvSsPP8gWf6kr+teUrDpBpDvQnegV4cy
W0+TLhiN1nn5nERT6TtQ+FspGtMfZzlGYeElEl6oWgMvlOehSaRSo5wwrlyP4RAU
ezbsZJU1/tSvz8TdCys6Xhau8Go7jRb9cpFk/VnrIZr8ju/hJ64i13CQPiAglcZR
p/dDcF5zFVvSRcicsz6WCZQhT4rxyCZv/VeM7LSV+C1MzEghYEd6+pI3laflzu6D
OLAOIxI7XhqDiVKPxIxyHR0K8UHnAZTc8K+hXvsqijk=
`pragma protect end_protected
