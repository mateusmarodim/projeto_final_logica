// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
T0l+fv4SxVM74/bkdz8yoI7EyJEL+erWct5J2A49TnvsI8PLGYMT/CCZUaPLO+xXFVC62ZPWZC4e
V0IA3e/Qgg1QPP+VdBnc8fKzMI4wXAA6bpiGBL5b8nFKr7wjt5hYkKM4r1H2ycJ0enu+oPJJtEBv
L1+4eFlXIA/g1UaMvpCc2ZbfUHnVJDfaBCxHTI7kna36M8QTT5i6uDb13v302yAmos4/+2v6nVMA
krZzwYazQZ/exophYY6g5ZiyQZEVec5xthPnn/8/KPaLI3FRIW0DDW4S7NqKzj9UhM8Wd9im2nQR
t9yULtFjj85VLgzivQYAlmXwELd6NFJmdprPVg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
TUEiZjPc4sQNm37FkuRs2Y4R/IYCoVQxeyhGOfZH4bE90gHc2IMEnhnLn7VCgCB/chJiNWb5PkRO
ViU9uFHmdcurQOXAWHvu1ip0TmJQKyxZNlCE8KmlXQggi9veP36RbQ6uZEH6oxQZ0LIRxiSlx0Pm
85jk7WdyGe4KJNsDeXQuJrR4T+1wku23GtL8DXrKIPcKpG0nXoT9fhmgOnLe9pOtkAaYHg3gGiSj
BZkTbDH1M57cqgKolvDCmqtDtTGp2CMfsGBfnsa0eOHM2yoQHI3DmQxK8h3kbO61aghBlGwFD3kB
rVye7wXehvoyE82fwKB9l/GszSBxHMSyiIZjRGL88CWDMRax8Tf7cd49AeCnC2xsSZwWK98almY9
MEn2i1PqBx0Apz77vl3RK6/rdUPd3jFkbZnFgt3qEZtYc46uOQ584OmNfhufTVr7mDpe9buvtmJc
6ADl8p7AbHtQRBjB+PeBuVvact1hvIbXcsIGkXGt29cXbwtPmKSAZU8s5FwPhujcmZ/A83E7eSX4
ZeDN2qivr6opB1gr5ILeh8wvZU2/D59PHVc1YsvTzcg2qjtznYdUEk672sxRLyI2X0cF/ES3TCi2
uPcHDhLDS71mCNmoKwEHWSDG0rZqVQtzOcXDDnvZ3XhlfRDI02k8ldwX5BK5MnL4eVFBpPBk9Fu9
2B6t6HwedOOVivXZ4d7DtDaJM5Cfq02zu2R6dSjAO9tex47pGXLXVxjK8SW1/aJt6O/lxX8MWzUq
WdFqD/580KD/cZKwwytiXX4+//l7et/vBvnsjproMo2f7c3WQbA0Cw2/Y2N8EjU3aBX47hNifASf
CzLbOeWo3eEVYg/jMjfVjqQzWQb+u1XDyY6CbgOOlT4Qf4QqJAgM6NKckA8uUMOi8e6U2aG8xgUh
i5LxwZNrPWV32niLVaPb7NP+TPCvvPvbmfwO6b0X1ASE+sHB/awMevJEVR/CMrPy5yYVFXF3QjCk
LiZHcbI20DFyu7omlpRtgAygtxlGvTQhMdENglSF2MdsYVXZPjfEIqAiMGvcgs+qRha0z2F+9eVC
bUkL4dfr8AsqcIqTiGFOM359BOmKkZahIUgh5s3rv3iYApAMaUdHcBd6cF/OEGJusNiJlOP7dEX5
KJcJgF16W2ncZZ/pgwnKnm/GaMoUCAgMl0ILV52/BNI4/9bcpfBxhly/aOLGhoJPIsKVr6zsbu+L
hu7r5sP5jJ9fQrsYmSsKpQf/7pL8R0WZaOCvJdU2ES6L6UXkwFtJFxH1J7Zp2AQo5H7u22LbtM8E
tIaRzO3EDOGMFFAtN1YtcyLu7Utk/OWGfmCyex1kBgLxTgPZgXqg5cuDJNZCKGjS6AtnMl0qu+jt
9OIrsHFH8wTajbqfR0V173pod+obbVOpLaI/1Fs4zQuiiBX2OtcgFqLwMdi9ghTk+f/S6x4c6naW
LFIMkKxU+sMy2YKeziX1aF++WMuY8C9kKwAdFaIpXQaYNL3wNl6UXrf6RjLlgXx3Q3bv1bVSkjvX
JAC3bisv7G/QFE11SBIPZZHCcNdtaljp1FFr6aPDNFYrMaSAoVVyyomzyzuIxXGgXULo7ccKtWPs
ZAPca+Ln3Q0YvNwU9H7QSJq1uDqGdkPH8IZuem/RWtG2qcrkv1d61j/UCD6C93XlDTahEtz3TQd5
RUhbC4uQ6nvCD+fga1BzDIVbN/eKCwVZpLM3cukyrNzBcZxwGjfXj8eDsDVEo5agRn42KRhji/Ua
bLh2E8rmjpNnQBeU0mxdjgLMj1eIB+P0jaBQilKz3qZYgvB4f6KJerg/U4b96zduZjmG6+kFf8ZD
g317mcU9BQQ7NSbeAPujbUnn//l7SNNeFbrOvsMak+L0YqXDNaoWc37qZeeiX/VLno6EZExXOyHf
+Xq32BYtb4qYuaT4icZ1Kw3zKjqed+dv6U50raRRINLgAiqTlA4DsicXQvaeQDMbtgvMfKjXzks8
uQQSM/e9TZjH0klG8MQSRXYB27aTdH9oNirGLBbzk7EeISUZQJGr2DRZFQjOEutKs6p7inrqNm+n
8Tl0BAETOxsKTZy+/zOffLCoGocLkxInRXKb7rHi9HYi66uKJnRw+RpxO6znKnb7E17XpMbm78rX
pleX2zS9AONoUlZjpiixbqIzG+VAhiaQUEkXP7fw3IFLX/cmNtrQ88+R3PSOTUcE6s4+hfbSbDzS
LUrts9nJvgqWDcABSXcG4H3QplyX8qDfvnls45G0KmuwskGCKypt8sTpQVn3o7B3TyhaqlixIrz2
XrhoogX3o2iEksoPB+Z0dN88iKwz6aANM1SztHHv4ndGtLPIwtHJ44Ao6jzuygl2/WS4GhHuhlrd
n7GAVg0mMHmXSuCek9slXXIlmgEk0BSVnsauGbleyNH8FPbDYsYHdWRktoPTASf0bgel0d1YRi80
68tWDavMRDbMWSNl8Zu/1CEHotLS+Xw0kTzKs8p7g8qUeEPQfTKAZgHOdBxOV9gpBc3BCp5iTdDY
sXHkygejyJ+3bsy9gQZOyaymvhk1DRYT53NKqdrNPRmA6X0OQBvYHwAEm8urzw1iSzMHoya2z1D6
gSwzl3l3Iq4JbXTKmtYsIpRbQf5MKloWvuhbBpRev6GvLz9qhDuBDqXl0KEosbg8XUZgSf8Vlfm1
UZnecmlXQkitnMTY5DYSb7LeiJLZDj1T/POTlskdiGry8+i2T9xd6wDy12JGdti73nVyjX1RpP3i
k1B1Qm/se1F4Nvs8IhTBPasvO5LcHvewcouaMxyYsHtTXtipsErd6iRDeMqWexlstcuCMcXWAOs9
pnGxeEdKLNgixA/ZBisNILwgBPOo3U8LBxMkCmToiWdXwSIECIDmxNo7gZUBU/yQCzs7JYGAHT++
edSOo9bpYNfBS4lxt+6Q1W76w/1x4YmQ18bmZdcZIsyT19uiZu6cltwOCM1zs0m2R9J4ULsdmClv
8bW/GSNvJeG53yckUFSlQ3ayFLyjl9C4xhrVKsGwb3FPnl9P52BXFnuyPKz+i5i127EaHk7rJ4YZ
iHwYyHXlobc7v86LBocFl0vlmYvBqspWONxW35UMgsoTjCfeeRGY/1xYv3jIG2QBpZ7mMIHvhy3z
ZlknL6CAwBLixkgDwYkc/OwjH5gZyEgou7+fHa15ybN/sfgw5Wmf6HPS/PCiqFi3txJWOmhTFxaT
nP4lREn7OUfCGKsRpBOZsaiWIkAXz1CGp2PShXSTYNDS+vOI+ZK6jIpFKIHC7XbieJBkwY3K1wNb
47CpdFSyW0wsmy+KZao2OteAzJzC6+iepPZyFMZXsiMmk2HerGWPPQXzuMsQI3FDWNIeJTu9/hX6
qLFgTjKb9g1WU4cgYYr0m6P5V46pOjs15ymh8H82owWdeQF4cCx6hgboBi+QnKlXkZ7Lx5J+83cN
T2b134CIpAiyGGaUnIo/z+r1irOClCP59fD9oSaUYV5jPIBsawrUghLqhg+e12kvmLLYoMtYaWPC
okS5Qb67FQZ1MbtVAghW+H7Vkng+bfpu6GjFCyDoTQtYlWAvseZhiOE1qx/YQiBaevDQjnUh5o0s
xC2KAG7SOoJ8J3KddWi8SSIT205qvFiFlHijEbXNMyks773darmOi3kq58GNoHw0bGjp5ShKdIA1
R0sVDpO0qn/eMEGr2fcaH7/Cv+6vd/NhoG5RkquY7Zr3WaRXGA6Ywo9dHkxp+9qfc8Qh+ZLKVH2P
HQvAHEPALIQCEJQi+TSzbp46xuprv1XYa7zGWERD4kOMujwvN32UT7rAdTlDp0PpwSQ0RnEUrbqZ
OAnqMlCfviLO9FSTBTCi5wpT5oGcWL6oSRRT6JKmr7mT4mA36D0gRjH4OHn2uPGRTikhoiH1B0WO
E1EfugJ2v1IWIujTZLT55QgeQ1dSyRxkAHBctn8779TLzKcMGyusJyVpUlYVkM4DI7QGAa1LhYkS
1UwLvzdgZOXKazqd98g//3yEFay2K2Rgygqfu6J0v0W6l8v83agyVum1KqHO3i/ZQCDkQTZH4B8X
qCAKqGylDmD8fbvNpqLtaYL9Gh7QOSlQDVbntz04A4ogNUH0IF9F2amk9tAgb095lDcWZE3MGC7z
H6Z6jApWlwMLoL3dJQBeVY1MgRve7qppae+UB05Q9O0i9TOxOmQ859zDVNSPM0QdkaIGHnCus+LG
5wGd27plU54O9AqphLat51ZMo9sMqcrR9yPX8D0WNY+MzIyVooGDjpt2WJzlqBRgiOFL7VtK2kkQ
WGxfllwVbHogMrDy+Iz71ujEnBRvnS9FXeVJj8Xmlbj4QrXw7xs4DhbSBb12HhzHZdrGoH56jAt7
5u0m/kRt/D75JOzbBcJOsTntilbBY/a39mNNSBC2gZZvapkEgS/BVInNQ88SW9ZanFqOSIPFo8AW
vVTYoALqaF+U/tWRI7bkhrr/bxKTGI5+BK5buYBl/atQI/2+klk6ymbpPFT8bgGMua9FSjKb2Htl
W3xYFaeSvULy9/dxO7mK3zOgyiyChdUVVoFVRAZiJScokcbfBtOCyS1IWPb9lXE+JpzzsWO6B56I
8/kFHU6gBbM57C1+gIrlD7bOtuTaGvQxgCfUdAwVBife6k1AGM9Sr2mUKu0ZtI6VA1D1xi47alu9
s1PmSfK70cd/UF/EjQvRaX03+l6m0sVO1QnLsWndzfMs1qq+UjL6hHkQUJCL+vOBImWqCTYNib12
8xGVyocPu/RkdN7sbTaK3HQAxIwrKnL3iE6IpAcHkXT0AUqFi9bWMn0pXnXRb3H3SBuVUagpGf2r
zFjmwrPffYUZ7NwZ4Y0+3ZxHD/BbGQ2GD0ezuJtAkBoHSKeuvcPFYzWeGGcq+611kz0v9muY/lCr
wrgf3hAO/oNvezGjWMPUmute6kZHmAHI3VE0cmfPkmr23FXocq80boWCXR8ctCjOP7YYcKav8v0t
5str/r56EzZadbb2goRCsQdVPvnNIUUX0oXMokER4H0+gFc5repMPu3ale+EDf7n/qW6EJEDKw6s
cHy4P519OQmFaDsyO9AMaJA4XnLTgTj40ezFS/UGglX6iokhXbKl2H3XaWVIPWYXzwCkQKD3zIMd
MyHlp3LhW4R9x/Taxt4Ikh+xcWanv5SECMQSyNhu6paWf8UY1KN5uxk9WZsQR3WsfKqA3wh6X0Xi
nc7GPadR69KS0QsRQ2F/3R0hu2X/JBlXvgOQh40/Yx7X58kB2r1rWH6O+AxyvvPV5R5jZPcJEZSZ
E0ecYwZNxtItfwsNQkKHdoJ+44rY4cYBPxhI/GkWWvpsV+of9zXPOo9oUubnS24ZskRoB+egup1g
zE5wJIHwQamVqn3YYQhGp2r1egh7IB2Wcnndj0Gp00onAm03jvmVR2jcgs7tK0y9NKp15N6YKK1A
xXsHcQzwpo3oRFFoPsyuSOj9nW621tOBCdzXoPDNRLDPVNUMU7iF7ZeZ9dHDVWIULwfR+hSGVnZN
4qxwQGmkl1n+i1043DWIUd31yHQfziKlMMf+dM5kUYCaI9cOz9vATHbHcTdruQN/aGUMHzkPL3mR
ckoIT4D9CvYNgCtplAxqPTjRkgv8H0OKRUZvKq4/Ug8VkYSzdtmaemdPbFUFn5SP7t6JOcNCXcul
GD5PCwY7ydZeVjUeDQDRDeDSDu6CkgW1iDBgGiDTRCTgDoPpSSrTlK5fyYRb1Odg7k/rlFLchxIh
4BRgvhXo09mleVpT4g5pZmx1+Ox14hpCKQoUGpigkWVpyobS3xsNzq13E16gISoXITl/NXIsoXv1
JRxtJ/fCgL98UvxzoIdzAY+MuooWFUnh5li/gLV4v04DT6wPcX5RWsqPvMSeSW2u7vM+QQj+EIeZ
/uwMh5yF/fhW3llbZbAQKIm8F2B/tigJOYFXRrSD1f46NHewUxDKGpSMPPcF4QxOqg9/J58mqD6R
I0aow3nxSAeBLeMdGa4WhVh+ajWPa7C8SAY9+eJ80/CfBqkT3jRy/xJw6yFSa7qzNAdwLGALq2ZH
2qpgGtW+pOeRNs+tD+al/5Lc+3HHLUsi1EOPmNJe8YZjqdxVxgWhCRvGRlesdp5dFw2bfNrv0F9b
/WhA6HquUnSE2aRCu/Q1UKkDiAsgphKq29Mn1wmtHX6V+2n4Y247dvTBFUl7VoT+bLqnbmIPMTXm
c4A5MHNivS8p4UCVDZk11xWeUaq+dxeerWOUC1KuPsUBa+kScptrmlloUQfXHex+HttAYdABIPSs
wSzBALJJDpxor7dfgio/EORR82vieJ41HloKeb5AoTwFly7kr6tmAYZqvJiseT2Vqp8KoRDVsBoh
c0u17c3l9iZeMaZDZbBzBEPWIWsD/WvdsE637WFv5iivSSjU9F2rVwhJTKcff0cMu9VGxUFCNSrH
713t0L7So3RLgpgvZQ8vXThIkaAD2lhxHvW9IH91Hq3vFYMVIQ+l2GDYhwjxNTNC0abLnl1J9dQL
g9TfzDEpOkd67I1hFQ2D2xb/Efx84ThUTwSOzWfjY+OyFU8/w4crH40vlZj0QUgtcTz/MZ8sOFx5
/1CF+SJGri7InZzhd9IlrSvb1ZZTxK/x8HRXayTZrWDVebGkxtEes73H2+tWpw8wNmF8qFFQvLd6
e+u/oTtyQ0F+lsrFwNEtMSiDKFdxMMHWiOrD5QaolTSfdABx4FKWiVCVFOrZGYQ7v/eadGFkdtHb
AXAFVL70Ol1BGIbLDBjRN2IeU8eiM4BwJ7NeC70qs8wimDRukHPtNVl0aJveYtF31VnkcmMzivzX
Je0B4e1CWDy4Ts4HGn2xQTYDNKG1qPM2MbetOGlzecdaQu/6xp/DJdhdE6tF7uF0V5t1IWIfDlOh
tEySQyAwjT0DgoNA6m6/250WBpGTDBxEYGnleR8uM0OYUdG9fiWoz5OZJKjaVsf32a8PBs89wIwt
9xWL5tUYSvnzaDlDlIcWWbb4yQ6GBpXZGFEr8ce8XqOlrZt8yeHh00P90b42xshHFsRbEFidJos4
u4htPdAbojmIB9MaV5CyHzNwMLCaQ3btevbUVStlONtb/JtiNk/MysJ3LOxRZX5wUR/D/QVF19ZD
uxQYrg5y9N+QsavNMe6W+XBai+ieCYlZuAld1Df/BwJd8UR8jIj6fdg5IxIV3B8N6uAdVvD97cif
2Qg5tOfN0m8tAeHi3onC73H2HtJlK9qeJnSno8oLQVCi2SiqDTv35uPq6YyZlYtbat27qinJyBWW
FbQk/1Q+V4N86SBie8xXVLQ6n1uz2/7aEMWyJJ1sc9gse/GbWRFExDON9Z+uQXrP3BCfEEOJ6l/E
wfjXt2ZFK7JZP9LtZCLJ3La4uvqC07tW8W71KbPIcOE2iSy2n9ITr2KfJVQ0plVaeSGCqvtOfQb+
jmCPH4h+k/QwFMKfkK9v1qhuRHNvtjjlo3fr91eX0oSCFi6Q2X4fqwOyo2BDCB3r7hWGexXViTt8
wFUWKaLD0pjNFOfy6dE6DKSIerwtKk2w1+FpGfYVMiVNIcpxO71/EdG4i/dVwg==
`pragma protect end_protected
