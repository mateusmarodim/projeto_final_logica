��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�:����ng�DSw]u`HР_��G���<6h���LV�laD=tp8F�C��*6�G�u�>��N5d�̬O�w;�vA���hgf��֛n��S���ڇ?vz�p��\��®g4�!X��%��2�\,h 	w�(  ����"��7�r�?���Ԓ摚L�U��x�5$l�eJ)�^p�޴�5������O$�)��,� O��l��<�*!?4�e���'����I"�-�ٗS��{���ِ�w�di��#�\�QDTF��������}z���χ�1R��PV��t~�X?��B��L�e/�!t:��N� ����4a��RJ��@Q�6�/����g��y@����wBJ^�qO�Z6Lˋ�<#�؅����}3?����/M���Y�
wp���6
ˑ�{�::n1���#e���!QK �aД�7n ��3�6��+��X�E��&:_m�	�jSj�Wq��>h������b��,�O��m�Se��0���)�f��ց~�k��>�$��D�O�c��#	���|b��,A~U��m�6F<9�jfM�4@�q�v�gv@C?i���[�t��6t����m!P��,�]�G�\�ʩt�H=�wK[���B��2O|*��
Dr�������=�[/|*T��s��Ec���l~��&.��^E����a��H.�$R6Sͭs�mK|�W:4�ς8X�"�c(`�c�U���)�I��b��c�R��=�37'��S���v"��4�:���f[)��g��\`��~��9_���am��;r]\�sa�������䑖R�,��6j�O�����p�,yZW�_�&�@yp+��U�9E1�V-����-���� b%��`Q��S�ʮL�YN���U�d��h���jNfi��U�ɡm���S�fމ��n�>뭀"/�&����a�ҔگYGj���P��Z��kVD���=p�$lD�f�-��șG���y��G�{ޮ���`QR�G	�	��g�׬Y��:C�1
.�v�Д�3��
�iN�� �:.�M����z�dC-�9�7> :���I��X΢|�fę+g�e�z]ܪ^����eWQs��>�)�-yv���~�y�-��"�����YBgMR�[�n*��!>�����	��+��N�q;��뭏<~ _�Tj�w�,Is�۔W]��[�PY�Ӡ�+�9\&�r����Ӳ|����g}<̋3 �ݏ�i���d�ˉ�)EyG8�����m�T�V��_C�s�wU��*#�e��}�u킟5D�I��NP�^�0�2�� ��g��F���%�R�-��̣4��eU7���EN z�e����t�O���(��-�L*��<��Ǎ;��ϔ�r�h�����s��|��U6�3]�]i0w�?%x�Y�z�'��1Y3�d,��);{�����^F�����3�`���e���2�����"`���A�$!���V���
aK��~"0�3b#�I�Br��/"(��ګ��6 s��ǆ��7Y.������J�������p�|��n���1��^U�r(�|��ĩ�*�m��&,<v�d���!�=.�wX*b6G�ϱܞ�o��H�u��%h��UT�kA���-�d%�!&�N(նƘ̊�*�W�ɻ�I|=�@>�]���(�[x��>�����_$�]�q����:�#6]��?�.�:�i�9���)i����Ev���TP��<V���E���s�f������ݼ{a�oT���)��(9��4��~�:�г~�v\�C ]-Q}�����
��s�xq	���?O�`(%�۞�H4���<{�pOe���CkOC7�)EjN0�!�|�C[����|�uX����|T_��9')���M)��D!�U��6�[��d������]N�����+�CJ�}��D����P�ϙ��bq�DC��dbZ��h�&����"���x	!��x�KUb��]��"�����c��x�p������J��ĳ�;<�e!�A�lV"1����D�����0~d��AYB%K�b��ب%*�)b-!eۙt�¹������A�a;�5����m}�_"(�/����Q3R/��z��&	�V���ZA/6R�{h����b����:�Xp�DE~�ċ6�N26��s,�g5}��Vۼ
wl;��ʟ7	c_����Y���c�V�7H����P]}���@��d؏ZH?�⪑E�-Ԣ��b������͹�6����������r�R���c��j+ſװz�Kz��]sn"���2x�Z:+,�p�;��HV,N�-���?��H*ΥrBwj�t���'��݋�,�2���!��hݥ&�N�A�ZMm���@�������YM�������Ņʀ-О�?�(��MQs�j����bHbAm��P�~j�ꜷ��x������� �gf
�C�J� �/�Z�B`�K�aA�`��������#Ñak{{#.���Y�O�0���Q`R�jtw�0lk�3{b�����ݔ>����"*R-� �T��\. ��5e��V�����O+����T�����#y~��y�б�?"��U��v	8Ձwh*��ůp���xj+��-�K������yl�=�!,�EZPh9YR��w���8#��J�ș�aJ~J���l�E�IA�Ab6�Q%����/�����M���~r*��^�.�B�3�z:- �N���^3�|q�@Y�	��ƿ�ܗ�z ��=���4�g��丘�xA�1�����W5n��]x��7��T�;���(�E��K�e' s�&�m�-QzAD�nWő��G?�J�����vL�`�~�o���n�N�W��*уeŪ^X��fKA�G��O��!)\Xuʃ��\:�z�Ky�mCeE/�p9~��Hy/�=jY��GbkF��kNbKԱV�$���9�YO1d�/��X�ic�Y����nxZ����2��Oo]�!�7WJu�z�d�;[`Єf8?�b@�غF�S�h��-R"c�g�Y0�잭��k�`j�l�GD�FɅ���]�L���4�:OF_�;�5ܺ�����6�Q�3�f0�+��б}�";�i��@a�y�!?ZC�6܎/��9�	 �<WW�|��q�/� ��P��A�$ЭZ���E�%� ����^����y��D��w�@���4A�u�͙��t���d�h�8�\�O�w�͗�vQq�B������h@b3�_˥��0ZC����)/�Փ�>�F��ɔ|%ڸz�� �SO�>�rj
L�p�����jIH	�CO�	�#K�Bˆmi�,1�G����]]��POtd?�=� 讜� ���9���2�B~�jF�bZ&Y��MVp�A���{�k���O5��y[���H`n����d~�k����=��G �A�2COF�9�_����A.J���w��#�n��]���v�)tsM��wc+�� K�02��p�����5����C�"�ҧF�;F�wF�LO�:�O���嶄�%X�r��S�t/��s#����p���B���آ�Ȱ��-]�Om��5/��o���D��C=L�O�hǬ���bG��O�F�H�E�U�_�{0�ޥ���_��,��e�/F�e�#'��D��7"2�)=e���6�W�J�h3���>������Ɛ�&��k���4�V�'<q l�*)4�6ޫ��9X�u �̰tS���k�;��*�@�p��lF��ݵ���8��IZ��b�+�(�LȐV�Nuå=BH�7\�	q�����?߇�� 6�=V:-���d6j!��";�
X[?�m��Vۭ֡]&�;�y�}��XO�'�'5O��gH]
T�Ow9��x	&����� Q�Tg���C3��F�����	E�!�Py�/�V{�9A���s�C-{BM�m%�y�cXz%/�j����\�m{�ɞا�cS�Hh�qk���-���m��W+A�6�a�1�j���k��h�*I?�Z�.��d�xL���%��=0�)m(��ȉ�瘜6<l"���,�o# �ܫ��L0υQ����RF~�LO)���VZ�]���z��mBШO��i��/|�)?�u�w��Н:ZV3"<ʞW��nاڙl����h�\�mH>�Y"m�/ݓ�����F���?h�ɓ{~��._0t����?�x�S���(��#GӚ�*t��X��Q���ByR�
�X�,_���X�4��!}/.A�N#���=�w;��ޖjQNl�8�AQ���)DA�5�Of`�l�cn��g$������$�UmL[���Y��iN
[-.Z���\�I䕵�ȿ,͖�PR�=6��&��.�5�.�"
�hO�q�F��ĩZ0���k��p� �Z�[�.��!��ib���`l���`5U��#�2�X
����
mu�r��9��B�Q&��QjOTt��pO�M��G�A�(�(Ŕ���޴�E`�,j}���O��L<	�b��=��8�OXzwQ��gU�-����R����m��1$*$�n�{xa��.A�s_�&1�� ��H� �E��&��GlL��M����j5"��`Tb/
�x�G�R����#"�iR�D8�J�����.@�a�J�Tq�*jQ�={�A�3�ږe�:ߔ�ǀ��uB[�z����?��4(� �޹�)%�3��9�o称/_���h�	���� ����
�lw�xV���D[W��� 6����@����}��'��P�pWp���/����q�Y�#?�4�(E���龷�6/��5��I� #���ԝD�_ϸf�`|UC|ǅ��)o&���D��h#�����&���ѻ^��$���~XڷFN_ �)���^��cw��@���nzw��R+rr �<��2�z��p�
0�S'�|� �wHc�ls�k��������X=���M�ݳ��h��h>Ά���\[��@~*{v���*�X+]=�8�+�m}6���1�K4si�ɑ�;�e'RҺ�X����[A��'�b�PN&����G���g{ß�	�b�.Mܳr��24���o��쌩`Si�@3uPZTdBӟ1���1!l�X�O���2vZ�0!��x-#��~�l&�9���Z����~4�{2x�0��ʵ��u#<�k��tU����h�ٍ9�.g���-�9��RD�\y�TVd
OC�� >�@vem��?�F��O�u&�N�
ra~(�8d�(��F��΍��x{K5�[跥,Q^��fhs{�z؜0��IW"�Rs��&���ZjZ�sr�K����L��i�u=�S�|E;｢��e9��$I%1�Cf����0l���WI��晤p��F�l^�s��^��y>��9�}[�Z��s����O��V�9 h2oz3ګaⓐ;�z��^������|`���8�E���ڊᰪ/R���Y.$��H��ɢ�ѕC���WF��Fa�;<y'�tq�E�����օ��`LY}�L����%�ߛ&�5@M��a+�B�͸��D�H��v���d�dh=�æD��@��xMTJ��m�5T����D�� 6@�{%_�+�F��b̦0-O� R�P�u<'�:�4G�� �h��Q	l~RH���
���)��W��&��E\��I<���1�t�i����궤��S��ؒ2��ћ/���X��mr�<$ʬQ;̐Y'J�*2v�m�X�:f��ə����nX�Il��I냬���Y\ki�+�,oq� �9�*]/s�+_=f��}ӱFv0�,����=�]�G|�r�I�I���}�?	L_���\[�ԥ�a�������f���uwg?��M� ��������x�A��?u^��cϐ�>ޝ�l^/�N���}����!�ٳ�M(�'����>���wp�(T�t%D(��~��W��ȥ .&)�`�ޕF8�sﮯ���4X�4�,��I�'�.���9�2�-�G|��"�y���#�aQל�FeI��s���8}��Zi;}��&��|��*+[���
{H�ҧ��ߠ;�O�(��1CU,���Я��?h�>��<F[3iAo�jf8'�6;Rh�l�O�i}C�%��'���Y�ʁ�y �sT�5#r�m���ɼ2�� o��a�[���?���n��{�IF�6r�6\��C�\��[��/�������fb��(�6��4��s�t8���-�v�ւL �th�L�����P���[�f��7��=���y�:9L��y2$!'����o+���$����/��{HO��<��"?��Μ*�s<����O�p-���m{Dr2̀�*�g�u�]�x��u'Kz��tR7��&ak��˝'X(��6_e�5*�.2'���,,��È|�<8У�[�9��17=�|��d�ZV���"n����: +2]n�+t��α�u�����W��.����6Ҹ�	~��IL/�&��k��N��#��5f ��9P�JX����EM�&ҡ[���
�?5&����=�n�[C��w��N;S��OpᲦ~虰#�͢Z�!��4hZ����6I�f��:���66���D��B��6����N0��5�I�����Օ��Ѕ���i7�<�`o��v̙(La�ֹ�϶���e©� �3�k�Ǉ�ۖ%�u��2���i��M?�V���>��x�>GV_��SieǛ{@�=��֖<Lo���%�=��	���KyHM�G�
�=p��9TP&>q/����6�vL#��4`9��D���)3+�`ր=Z	���Y��Z�CF�vP>�[��TK��o��� h���7Wp4���Tf��3ֶ���ߐ	�Ա����)���6yR����ƢΌ���������s֫�R�K��%i�c���M��J�O�2Ԁ���V?�}�oC�l�C���Mah����w��4�=��<b/������:DN�\�r�**"���t���~�/eۋ=� �'�$ ܷ0<	He=������0>��T ,�}Z>b!���KMg]���r��	��i����h�ql�Rm'�l7�﫛��\9a1#�6L�w��^Wc_��,�uR���[t�بƶ���`u} G�q�(%#�Ni�Mn���)sס���0�6�9�����S����1��H�����DT��w*�eĠ�Z�/R�
��#'�	����޲�7m):G��°@D����H�[ӎ�G�9�L)��	'W��E�	o8��p�r�x��y���Z�0ȗ���be��.�p���F�$ʹ�w��1:�*���q�G��Tw44c)���Y _^��9��� ��W4�/��K�L�F�+�ڐQ�n;Bg(�ɃQ���9���h��U�geu?e,Qp�qє�v*�h�$\Y>�u9�Y���T�֡��A��7�녻�>օg���U��+�՝J��w�at��}^���`6I�A\�-�h��{׻���z������C���£�t�H��~��{�r���3���'��B&�&"��]�q�p�9~r�1���9 O�`i�1�ٹ�P�x�[�(sO'�[�2�T6�~6e�gN��-.���q�G~���o��F,���Z[��U����,�VI�}��xt��?3Q4��<\��0�$�"���,9(pV&*�[r��"���HX�`^�7�����1|.��N��o��?	z�ar��}�F���2�j�&ś�`d�q:HlE4 n�0� �!lҴf���0�6�,v�� ���,����aNt�Q��0:���N�YV
1rݔ��P?D�`&�qIv0!>(�LE�=���-CP����Q7!�{������٦�a�6a2	�b��f�����`�z_��a�)FU��#���a\�]���I�=�/
h	�pakʦ�*y��d#x��?s�Tq�&�l;5n����O����
f���r�o�4���ȿ��)L����3yJ��U�p�|��+�v-e��W:�V���v4ca�8vY�C���b���0�������b^$}'�u�j��qe�:�D/q�r����k�$�h24��fE !�[ܡ3��i�����z�0S8Qs�:�hD�9���Is��=,I)��\,�O����G��Ɓź7+�o*���������^��9X��:̿	z͗�XS�.H�8G�x���I~������<~4�.ʠG��eg��
5�r�Y��8�ue�,�kz�����
i?�4�䶣��R�"�\��X��8�$�ɠ��y.e6lg
E �-E��W#�t%���v���J���'0�h;zn��d0�bVc�0Zd	4�]�j~9����1KJU�Մ<��"���UG��|"�h�GEշ��j0�g��F����.�q�K�LxB���jEKPO�%�j���j� �*�5��U�i���>r�*�vv�Ĕ�#,t,�a���n�V����z{�EN�M(�]�p�#O	����W�=�T�l�+@(7yU�p��@Yo��4ӵ���]Gd�l�����t>�ԏ	��(�P�4N3�r0�;Hwr	���R�wD����i/u?���ȣ�\�`B���]DS�d�,33�U�|u3B�~��� n,��j%�+��L��+�ɵ��n���b���3�V��Լ���t���t���" OI�B�=�,~����5��eo	�e��n9-���%{>&�o��&�[@�\Iw8d�'��8j#��y�\�u�"X+�|_��׉Qw%���y7{�	4H(��ʦo�4�"�˨v��^��OŲ޳*Ӟ�q�״l�����kF��Mhܬ]�r$�I.�鈠�hN��8�b������E%�㋎�����9}
d�1^��nj`���Jp8V!j/���R^R�,V��r��B0�7�Q ���[�������b��@[_��w�t�4
�ɋ�|�b��מ��(G��������k_b}$B_�(��
q#�l�ST$��8�<�r�E�e�X��(5I�W�n쵵i#?��v�j�_Ĝ�A{��S.,��wP���M {c�,0��Bb��A?������=���$��L�p����ڗ�_a��0µRe�
��Ȗ���"[�mߓ���E�S.���t�`��Kɧw.Ր!�i� x�3⽮?fo),f^c��'�C��H�qu�z�y�<�vi-]ݹ�Z�]���LH�f��<��ߚ���	b�ܐ�u�䴑H���	�.���	�+7��M,�>�
,+��'�R �HLL�݉`� L�1&3�
s�L��|�e,(�����v�i/���.�i}5QT����-}�����z�	��m����ǂ���e��Ҏ`v*!_���I�?�,�x�M���S���Bb�b��n*��/N1���M������ܝ�� b���Vlޕ���!<��.���M(������t��CBQ �7���k�"zax�E����\���� R?.�<s��9��1;�����b bB��_剈{Kn��H��K��\��c������A��K4��+!�uC�k�]�ũ��ւ~�3h_����Q)1M��P�,���z`���'I����8��7�EɯNr�� #Oc��\�i�ut;4�{��r+3��(�v�єU����I_ڡR����	6p�y�B��롓Y=f���ԠJ��.~���S��HV
�g&��h��>\���� vh����T�{�箹���	�������nw�N
�Kʹ�����IP���̠(�PjH�zlb����\��|��`f��$��� �%�Z����Ƒ��b"�.z��l�F1 �� s�����ҵ�B���� ����x"����N�[ ��u��!�C� �ϓ����}�FJ��,�G�n9y���UoW,��0(�|h��\�L'�+2����֝��������goHn/HW�쎾:�1�]����5� �CS��Ҡ��U��5Fg��U��<�^��-]�Y���r]�"��b=L�G�f_������`��&d�-0����w	�0~)(�ɓa]�CI&;)��J�4���ލ�V<�G�S���t�̞�C��8��d
�#�w��Bl��84��|����9׀|~v�j)�_ch]����ƻ�!�|!E��Y˶KL)�|%Tk����?�?��V�u�!�4���H<k�����K�Ҳ	��?%��GƵ�3��'|*l+��-����~�((���ς�"��|�G��=���{�����f���Hg�$?MV�M/r��|��;9�8�M�I"s&�lcu:#����4x��
^*��o�M�l��]�d�b.�٣dfo=�1F��l�9cyчk��,�y��H�����W�!�{C=�?�P3Y]E���z���s��h����͡Kb�������X�� z7��H'�e��"�R���俓��~[P�7^�"3�iTg�`����=82wj��n/*�7{^;���|�p":��L��#p�B��2|~�ɋ�^���-ʹ���l���3&`{*��X.�W��ҽ��B��Q�@�9��+�k0{�@M���/�O��-R���:n�������˨�T��� ��)s=�_hG��XrȋL�P�Bq�(C����.]�J�`$n��ɓ/��ڶ
�^$(�q�ϊn\�;�ն���on�Q8�~1p����ZR�Wp�J\���N탱.�7���s����Ǿu��q
,�홇������� �$.�<X4��k��?��nv���`�es���F�aH�D�G���I�?�0����:�&X��
-Z|>�^ˈZ�:����MN��\N :�%�ͩ�p2�k�kjE�U�=�n��hE�Z�c���z�m52��WH]eA��L�Y���fP��^N��� ����z�	�ȃ�@��%I��Zi`�1}H�����:�2���_6���s����|�A��93�D���75b�}|�Bڢ����b�����̹ǘ�Ek�e@���]r��:����Zxb�{�fOW�����hZ�8lY����zᕍˑ�?�m������{�m�Q��<w*V>�M����5 ��HYut��D��Ԙ�n�jE�������sf���s ��fށ�KT8%��P҇`JPX����	*�<��(P�G�^4���86�ڛ��0,آ�oy테��.���߷����$+�e�����r��\B�]@4����@�ݪ���ɕ�<#[�>C�n���g�V�,i��E�bS��e��0}\:n9*2��4:
�b�$��N�b������Y#���@��7]!�P���k�Һ�1'N�!�T�:��Xj'(F ձ�ت�ς�1��l��f�1��o:�,����j	���]|��'��3���17����q[���{��}s���|����BF�P����8�eG�tl�����s�pW�"�7{�[�������a}'m�|'\|�{��B#�Ԋ�Z����}o:X�"�2
��G+	��(���9
bF��⦍u����랊���>W��60���'��<T'��E�t�k?.kC��}��&$�kO�v��=�Jes=g�}
�������Ƨ5��7s�i�����!��ǵ�+�2��f�|e�%�dɾL����������23�fc<��{8����L�y�MU�X�+zV�N�O-bi��tH3��Ҫ!�����0�>���?j,���?A��ܶ�Y��uib� X�?s�brژ"�Oj_�I�t���y^[e\G�S[�����{��4��M����J�v� �ߣ�-����7�dy��C�>��N�N��(w�>�j���4��+a╀���&=�P����5��!�D�Ʈ��+�z9d�*9�R�yPrt�&3x)t&�V���;����n`h��A�b�#�����C��c�V�L��Й�_�|j4�z��5v�UT0����Y���_�K����.?��5�d��|k�T����AP�T#��@c[��#D�F�'v�-b��s�
�40��OL�(w�m��g�IUu'�{^���Zb9�X>��fm��)�+��}5���Xx�0��&^ZM���m��b)?HV|�����-�}W�"���mD@�� �ImEB� A(�1��*!�iY�`[٩E�{�1���Rsf}��ͺSd�؁sE��Y���K0���l.bՋa�`�1���w�`>uFțw��8��'�v�¯14��Q����IU�'"���r�l��F���x��a��;�U^ˆRr��y�a=�P�X�n���rv�M����'�]DgsVn��Z*�W�.�\NW� ��K���ad�UU��މ\|d�c��57Gٮ��l]��>��;��ĵ@�Y�4���D�N@)$�5�
(��M�\� ���N�]b_�$�@�$x��`��MZ��QA�S�����U߫��M�gÈ���0#K���Fץ��N�2����ߧ���ۘZa���শ�ng�U��T�,s�/��L������4��föp��J���d�K��^�P��4cNՌ�~��#�_e�i�̋� k6���WsD�:�K��H��l-lr�[,����~��B�Y������ݎ�QՅ���p��6��=��0��|��SY����C��go��^	�V�"&���/y�8W%�{��F�I�=�d"�9��?J��2e��[1۬
?F��� FQ�	 ��" �D3�Nr�A^���$���^�*_�H��I-'�k��ߥi���KQ�%��3�Z�8Ah���F4��#�<6���6�;�?*��HT=9(�ÀG���1�����)�T��w��8�B���L$i�w�vաx3'�S{���h @5�=�M�TqӑL�"����P{�UHƏZ�Z>w)�R���J> G`�2��~?d{��Ұb^`������$N�+��R��/�Q1h����_�js|JvaY��6u'-�1��&2���QH�'n���
�\�k�/���w�+w�D��f�9�[#��,��B�Z�Κ�������u����@��ˁ������?�����bZ|�(�̹���2��aʖ<�`wɹ/W��S�F��Z�k��w3�$������}�n�L�*�~ ��/-z���n�|��8q���o���+7mm���w�K���VA�/y�������:�t�x��K*2���y���B4���gmY!����&9L�/�`v���7UA�c\@�M�w{ڍ]1��XA`u��q�)�����d0��an�"��'���w.�/�1r�Ɍ����LZo�G�Ox���B�s1���?(��Z���T
�R���I��Q�qt�l ��N,)���Vo������U?�K�^�9��ok��}��塿�����B��>{X0��C��K:s�v����v�@ϟ�3I���K�
˘�"�n="V-q�c��،�� ^.M`���q�'&�s=j;w��6��=�#ӠǭՍ;��4K#�=|��� ��"jrL�~ϧ��[I$�Q��7�5��=`cPb��ð"saQ�-���C؁����Jjs�\F��_�n�	.`�-o1(��	SR@�PB��Eʑn�ps!P�{H%O}"jK��
�>�r���������n����H-�=u�.��Jqi�m.��	���b.���U(-yȴ��%��E��_]��I�7"5�! �[�T���\�J�MD�[��� �D&���18���1,:��Z�^�}cc�:���X�:��~���6�F7�|�#�<��1t���M?��J�Cq�d������&xy�${�Ll�>�n��������5�EF�v�	R>��eWOU�O�bb½ �op�;,�k���	%M�&�43���a����_`���	��D�ψXE7A��]��J�*Eڴ��wq8�?v/G���o�v!��	�p�7B2Lr�`�ߴ*���Ē�<�^v�c�P�q	�蛟j��)?�?��+���C�?;�70Q�-�¶C�fq7����D\6��,���p���1B���]D�)����nS�^+7z('X䨰uA[Ƨ@PR��|�$��Kov���Aqj:�L�]�n=���\6��d�{�ǆV1�E�8�����v��j��PWu7��	���!i�w�@[���W�H�W���L�]�ԍQ�~4��t�(�\��'�7��k��67��h��
�š�*��9#��F�V�3-�3��ɇ�>g�� �@<]ޘ�R���6Cy�d������$�WSZ�x;���:H%�Um2:�v��R�`M~d2گ�.FN�8E��D�1�R�ؒJS;0���8��/w�h.S����w��������_���~0��`�n�Qb��&���
��� ��=��Z��r�6�e��>�K�h�,�s��眒�i"��̸
�Gp�Ѻ���_ͤ6��C��� �Y���2��������Mɧ}K̷��a�<��ZrGq�'G��(7!�v���N3��}��9
W���"_��7�K+�o8�����@��s�-jn}�Ag&,�ɢ�8�����J�C�s�U���h7�T�C���\�Q]�]��e�x�A0�X���o-f�+2ی]Nk~A��Uc��12�r.^U����#_A
�>ٸ�A�B*��^gEmF�Ѣ(��t��������QPiִ�U�)�'�:�Ӧ��#�&_ w&ty	IL5���"VfXX(����ς��yE���AA��%��fյK�,7���S�ꃰ�$am(���f7�yO�@"XO����i�FVZ@(�琉�1�g[F���}�_|u&$`x�1fë���X�6�|zW�F��I[?��dL.]��-����.�H��=^��@̀����,��
��pR���nS�4���m4���#Y�]T���B���5�a���Y���9&(о+\�P&��'
% ]�=� g���4qxIA��Υ�h.�˗8�59m�����8����t�������*����}5��}*0㹲�9+Ӕ���OVe#����&s9�9��+N�;��6n���x,����> p��G3�YBJ;i��?6���	j4HZ4|we�hԼ]Cr�Qo���|��� �5�O��{<��6i.�l'�O(~�4�)a�=Y["�y#UC�9x�D�)L ��d�X��f��3r��dz�hk�J�dݝ��bkk���۴��-�V���Ƴ��݆J5�Χ������1!3{tRzH^#KV���ýWq"O8���<d��9��c�6���3I���a��[�l�j�wV��"���V0
��M�A��cQ�P@�`�w��r��;����㘠/�����Pkal�~�����b���Z���@��ˈe��e�\{f�Q��9gb�[���B���mϩqbٳ�E������� ��f���(o/DCCBܓ�ۗ(����\�3�ܕ�qPQ�f��$J`D����~5��}h��ߨ2�H�,z�������d�:GUQ3�����|a����N0wy��0����{�������^1B�۩r�>��ܭ4zo�n�7�h��CeLw�w
}h���m���Oʲpe��	������:&{=��Q��MO:͖YֻD�31e=��L���Q�q�_��d�6�}|�o�x�N�mM/Z޺����I˝����$N��T��d^ͫ�Q;�;��P_,W�"�:-E&���f~�����IZ�Lأ�~H�O�Y��A�]g���eT��6ov��-޺���:E��܁��WTv����2�0�>� TǦ�"˫��eQ>�(^5U�Sm0&��.�[�b�@��q�gl�]W���I�>�M���z�)�6Ũ�Lk� ��?��nD�@�=X!�m<H�l�y�܃ݮ��@�ڂT�|���H�����36O�C�`�kG�m뗖�!��O�I96��䷻F:hX�M��NM�g�1�<C3����C���b���k4��<�_˲�7�풵*%Q�$.-�x=���q���*<S���b1���y%YE
����k��'�T�̕EReS�^{�Q3���2���,�̃��}|
���S7f����v���$-/ Fxy�z�aڬG���F�B�bHt�R�
Ĺ�!��g�)��6@t�C��w�nk>Q�g�48m_|^�7F!MY�{�p�R��0�����W#.W9
�,���p��@��;�e�֚�nZ��u���[![�K|<�N|����O8���6~نY( (���^�j�6�F}�����?�U��Q�K�N��B��ekG�R����o���T^��j��:��I](����=�dXfD�ܜ�a��t�?�kG�װ�~$��ޔD�M�d�кZ��m}�!���P5�/�������#ȫ����Y��d�˻$� �=e�Ibݸ_J��Jf������^ 2�,P�>����V�yx�c-f�~6�0;=րR�S��m'�˩K���ܫ���1��K9�m3��E�F��j���<0�;V�}�Z"i�
ō���������zELN!3���A��p�ܟ��:�L"��e/���	�����E�gS�֟"C��I������O��x���j�����q���Bp�B;}uր�����ٿ��(zF��:�ԊE��2��"�s�HD��M�">9)E�P���ϑkO��ķ��bdy4����& �"�5��],���@�y��V�h��k�RKj�<rvP=M}�+�{__	�zת�tvf�|.� �?[&eA�N���3�J#��a��k�ur�����.�J}9���C�U�nߘ5'�*�8͗�{΢�N��Ң�=Ks�i4ϫ��֖uP�©	ixmY}�o��/o6����_�[��B~h�#�H��q���,����̓�j�Ή�|����[%��=^JQ��)Rz����ֈA�&S���>����It�Y��Е�W�&�,�(ݷb}�1m$��-I��Fw L�s`(AJ��`����m�Q}�{��5�C�ha� �^���!��v�Y8�4O&��ú[phk?�+&G�_|�Q��c9���6�o��?1w���,�\r���ޢ�OuJ|�S�wd���:�Q	�5�ߜZ���qtV4��,�)`Bҭģ�2�$ݠ^�NݽO�$�CU2[P[FSؒ�Kչq��!g�g`:p��!*�{�PѪ��6��/c����G�\�h��I���n:ys��]�%����GX�kўi��3���/�j�CfĂ���6{7ā�+�A�b[�$��\�n3�5�n���Z �F�^�E]�B�>�?"�q8[��!��e�y8@C'�-LӚ���l���SЉWX5-@�r��,3C�Rn�S��Nˋ�r�z��G�u�@q����񊢄���}��6�ɾ@-_�$�[�$q�* ����݈D:8� B�+h?�#�6_���e�>IV8�p��� 7M�B,r߼a1�9���JV�Q�.6�d{�y�9&~�	�R>!���Wj�e��Ư�N�}au���*�M�=m$O�F�]}m*����^J��pa,�\�"��"���썹*�U,ͬv���'M��RL��y���U�k�U������3��L#�8ܔ�2���)3���ՌH���,Iə��@����yb{�J9�>7Su��pl
Ud� Q$.Xx�l�_�l���ғ(is<���-�D��4;Q�3��W��y�nP}�lN�u).ooF6%Ԋ���C
J.�.�k��B�����3���(F"�؎����E�np�_��"
\�~g���VQ��$�>�$'c�"@����uh�g��N_�8*�{;���{�|�y��Ź����G���f���fr/EI���"]K
1܍ײ�,��?��&�W
CbN$��)C�?�?l��=���� �W{�I�iоepI���@�-A�;�~ �[{��得Ɵ�S�:<��:`$���x�M�vQ)<$����.�{4p�6�P����Q|��g�Q�l��/�d?��;L`g���w�5=�y@D��%��"�K��N�"�sx��8m����!,�m-�n{�%���cΚ�"���RA�,z9�u%�%��5���e����Q[w]K.Ij��J�5Nu��V_�붧Q��2�zo*Tiq]�^�����7:��7�q���۬���P��� ��ʺ.���#�����A�2Q�F:��Bh�l۩U�i���=��.R��G��{X��)0�O��r�K�S��=�as�	C~g�5qT�sl뼬��	(����x�qЕ��B��x���q's[��;5�%X�&!
h/n~���K�x�v��t�.'ک����7�����7<<0;	�~\���*�Gb�a>�����wii0��*��������q=���6eL���_�@�@m_̹�^�G�`�z����\	�?$_���H,�.l�����r5��{_��,���٨Uc�� e\;T����JN-�;ش����z�F� >�=���	qI?ֿ�������/�=�w�&k�AQk����<���%gt\@j�܁'�`r��Z:��`qZ%�t�����\s݉����ba7(Dj�Ӑ���bl����Pӯ��V����w��v���G�/(���MI[R����=���i%9z��(}.p�{�n� EzZ$wI���d�(��(9��M��G��I $�9	v�קEz��������<s�G�u�ӈ>m��e�i�yO�+�)�l�ЍW!]TJG����!�X�a	��~�$W�u��-`��(�Z0w�k;��̃������H����(��:՝W�Cîz4��&�u�k@�]W@d��ӆ�>��o*��+����^�`q�GG�o%���u��I��\��U�:�_q���u��@g%ԂI��Ϫ;M����*�Vč	��l%��,�n�����>�w5�#�@��'��N�W��]vd �I��6�K��]��qO�W�@���}T7�Xޥ�$��M�8f�=ȝ��=,�Խ�.��>+�#����ƂX2��xbo�j�� >�_�*Zw9b�n*� Ue�k�@������@y��d�Ib�Z,���a~\@�E�#{�5����˞]�enu��H��s��c�O=^j���t�A��:�l�Mc..��K��t�z��D.S��X��3*C�Ǘ��|C^)~�������jO!Ƿ%�h;�=�",�h���`��:�!�cO��!MQ���aA#V6�?�����^�K9	�zQ�S�7�I�P�q�&6uܒ��������%�X��PО!��wk]1�<�!�|���p)��/AdO����
�X�Zeϧ M�v������ !�T��ǽ66X�W�*��JX�p�;@���ڧ��i*�W��y�i�Q�:8Г-�3��?`L�^�h��GU��pD��嬗|�T
�����<u<�e�� g���V7>��8hƬ��$��ꏜnm��TB7�uc ꠑ�&���N�КS�J�[��f�:YT}��sf ���\�Z��bz1Ii�'kf��/�a ����m0B�e&)CjVX3��04�
R��QC�v	�ۭI�W�������I��9��z���כ����I#��P��P���S��W��@0��4=��1H���;�!��d���:D�K#S��Q��e�7�%`iaJf�r�F)CX�e�ߐ>�'G�{��g�����2�,���}��]=�����x�N�G�g@�	��+�b��o�(7�Jƙ��q^&s�2I�d����<	g�]e|vCyw��;Z��s�h�r�Z@��Z�a������(&d�L h�#�G�0�(.A����:�t����6o+(�����n��*d`��;��|�x�B�t�3
���|xץ�܇$�` c����#�Qiܸc{��t����IS?��`����w]Y����NL�7e�f�A�Ip8ml�lE���
\����i�v�w�-PqbF1Rz�WQ���l�Wx�El(A��g��@�U{Bt����Az��m;�����v��nߏ�U��X���ڃ�oԇ�.�k���4c���!:)�>�IpE���ы�����oK�uf.57��%�|�;��A����Dn��#�Y�-���:��+z�]�ma�'P�\@�۵"�.��b���WtP|
Q<�m�0ABi���P��$�l+���[$�c��XA��u.�G��8j|:�Lw��³�&���:�k�Gqt��,c����*�r�����D*<�G}�ï��=#�F��Y�,��1G���8p��n�ۗ[��Z|eo<M��z[����\���*��ԃnu�| ?Ę�8��#Ux����/��Q��[�3\yا�)��
�f�ƻ�����Xͣ��q-]s�-'����K�#2�V��7u��ӟĉ\ւ�����r�ys�b�j�j��hb!ٿ�P�p/v�q0�`a��*É�ѿ�#�\���U��*>X$��(��-���¦��mhe-�cN��2����D��X័�>v�a�O�ː��/��)�{��0"J5�nۣ0)����,/i�ZUF�ލW�p<]�'�'��
���_c�Q��*�m ����@�8������i�B;��M�A��!b�WC[��{�懑j����U�ӗ;�� l� ��WWF!]G�������?y(+�����������B� K�|;�Y�)l�	`[������2�%P�b���'��@�Ԃ?��(�%rQ�$P��e�l\"�3�rø����&�����2�[�b�K_�fFܒ���K�i���v�/�7��-e��8;�3�n��n�������f�[�/{���j�%E�� �1�Cl�3�U��å�u�p��1a:Y�q� 0�����.�2�zzPWe
8�9�13�;Hms�3����c��F��sƣ�ƿ�!j.|��u��Gi^d�x�w��Z�DR��x�{��?�;���Y4�$�P�%�8xvF���������iZ<�� :�ڿ��h�m�yN�ݶ�D�����z��mA��&v=��� �����d8�˷��cvVL[�2��[�.��yJK >9���������z5
�%�uK�K�υ7/���RN_��>�1)Э:�5 o2�����������}a�H��m���ֆ���x0%��l+:_�p�/�F�e��M�
dw����H���%2b�H��F�hd�����P4@R���)e�K,?1F�,�@��`����w��&�>fE�׀�:�>s=���b��J�X�f)���>��?�	�ZB;���;�61����x�zk�
� �+��HOn�%
��"�C#"xv�}�r>B~E�W�G�$�/�.��Ofy��p%3�]��ݮ��@󀥷��?�<m:���"lͥ�
�RQ���0Jar,!��t��zܤ���5�؜B�6��@P=*^�y��X �l�(~;.�f��V����U�l%�M�'��T#��Fix9��Md	��)C��s�� R��� �rUZ�ߴ�v�'ߦ}d֯�g�Ț�p�
��&m��.H���2�&t�p
��Eq8����|��d@�͵����x^�����	���މ�$��)|4l>Cn�Fӕ�!�#�)�Q_�p��6���'�V��%%��D�cג{K,��74�'��22��eʼp��j1��^��L����+Z���Z��D�\as�T��nv�\���@�EW�|�o��z�n*7���ʬ`�"|Z�g��jkk����^��!�}��:���s��Mj���`!��4����_�U�<O����q<�{�U�4�(&��fb�P^���
��FR���!T��˶�r�M��Q�>����<t�Uv�V̘'�W��X�6�cC|�?߾G9������ȤV�[�2J�4�����B������yZ\{���>Ø��u�@�������	�ک���P��"�4,?������=1lp��򫱘ֻ��W6Q�My�F$���p_�z���Ӡ���]�_0���	����$��-\/n��p�ș��v�Y����m�S%t�-�jh�|�]��0*|d�%4$k��϶�k�����W.�{0��c.;6�*}qd%D��,�ޮ�ks ��Q;�Crǉ�>mUb�[N���ȅ�L0/�û�/�=j��.Fq���%�y�T�r�uU���u?1n��c[�ϧ��#�Q�F&�D&��o���[��e�،{欎k���{�}��m��ю="︒F�܄4��`�$��tH����?͓�ڏ�M��Nd���!�i.�D�E�N�'嵁���Lv�V��ЋD%��(����t0߂�Ƌ��ښ5kvZ��Zv%}��<��ˍ��s����C�Pb�ʕ�q��g�LS�dy�a�kUޞ��-�O�Ll�/�]Vi����� ��1�$�F}��ϼ�x�:�׺F�/fɶ��b���\��僺���_��`B)���k�+�&��A���Mwq�1lq,�Xtn����\�I�<��x"cCJ;Y�
�a�n��á˓�.bBviD&�qa�_�NN���#M>�J�����P�i-p**/�N�k~2`�������� �-_{BmZ�$Yb�$lJ"@�YC�/E��m�� A2o8����go�憛����k���R�rU�Y>eIӖ:�*?�E�����xI)����b�>��/��k�Q��VYT�w�1��hi'�o�u$ ��*kxm�y5)^��O�@\������#��@:	6, α��	�,RO�Y��٠��7����:��K�ς�wf��M�V�[_�V���������K����&�����K�s 
Eb�|r�m�t ��(�čeQ?Ԣ�8����g�,����c>�~>�<�jJ�`c!�FKL��b�a�^��|�[�h�{6�&��lՋ�p�]���[fˠ˪�����X?r�7N\��#��Z`��x�[��^�-��!l]��G�/3�б{�$T'T�*��%�c�E�����S�4,��������7��e&�.G�al�d�U��g�F�!�B�YyWg׋XrDDW3�M���z���z^�cJ�hO����W-^�@���T���6)���,6�&�Gs�n�1m�K	ь7�h��ʁ��ۑ@K՛�S�-	�;9�q(�hk�"o�+�����G�%R�g�2�XF�:(�|F��@(���f_����O)Ez������4��T�q�=���:�bc֯�7f0��н]�p#��_�)aYQe<x��Yz����SqJR�{���>�WY�1�Po��:����W����U���,���/P_i��0�cv�ea&?���m%�������(.Z�74>h�:�D�GoM ��U8V��f��d\DՕ�F�sҗW}p�?hG�m!�;&�Y�TN�;�����Ra���A&zR��(�X4��l���Io֊Y���y������9����KӴ9v�-~�2���P���ޏ�<C������0 ��J�h$�s��L_V�Z��1D���{ Z#(�O��JW���<�9��;��\/�|��@,�R�soa.��)&����^I�4�K!��F՛ʤg�(�V~��)M�q3�]2��U��s����Q\�8*���97�����x,�J�:���*�&��3�v�gD\�M�� &.�t�9��Ѡ����E��b�T�ߴ�e��\dzڧkR9�죐����2D�|غ*�@��4fJæ�*5u�J*U���H�k�3�լ_�
D����Ϧ��ʆk�\5P��zz�)8��ɇX�@~���F�OD�wa�l�y\^{���5�M��57kG��<u����Ne���a�����H����H�	5�NV8�C�ض�����ТT6If\��O��Ʀ(�Q �ku��y��C�bX�:<�},S��(L��V�Ðr7�8�`��<�ǲZ�Z���TK�@ߩg篎����KnV��q���Y��<�#9`⩢���L�W��Y�,��&GP�$���3�Z��C2+����r�YX��k��`v���f�S>�ݖ�qػ�s˖:�����|#���<ҕ�/�����΢�+N<ώ��͠�]{�n����Ǐ�.������ 8a����h�0l=�2�z��s�S�g��g����n��)B}���$f�L�tu�W.F�`���~�D@����{�j�7�!�Jd�ѳD�L#{h�^���I;-{���ši�d5�}� |��0����;y��U��NeO�[S�#6�A���5Pv��<�<E~=�ax�'?Ti����d	��x�C�|�.�)#���"���ьO�?����N-�(��wv3�1HWcN�{���������)�b���tE1�fa��Gl9�M���x�6ح:hCOC��]x8�P��FyJ�B�B���l����KQ���rB3Ǣ��v!���@'����毙B�y_���h�`r^���/0��qs��"�'+�]�q_,�b���"���h;���%��=�Ás����t94=)��崹�|z���͐����.�>��	;�K����Ĭ�Ῥs%� 5�½S]��;L�PV0֓�䔔�r��}S&��V5D�\&���y��Z���ŋ�H,��\�t跶'�������)d�F�q������~�,���7\�<�PC�p@�ێ�`*~�gU���Ws�(h�o�N�6i`=SΖ>eק���V�Ί�E�y����Ǯ)�o&>du����E�3v�4|4h�J=�+N�r�E�*�e�@�(.63�+�6Y�w.�sBT�O�+�3���{��i(0P$��Ȕ�qץ�Mɭ؜�#逍}I����W��ݔ�E5�L�E*�P�a������GSȽ#�B�R���S��ۛ�
6`9Dmun 8p
ڻ�y��{��!h��}��D��SZ�2^գi�؎r;#�(xN�L@?$�d��l�Q����Ï�`�����͕�����m����Cѕ̙V�����|�I5h���l��$�7�<4�NJ4ȿ���J����ђ2�#�6�d�-�A����H�;����S��6��T�w-D|'�^���\�D3-��8`^q��������s��0����I�k5��Rpw�ȿ��"���|����>����{�.3}8	��H��n_f�Tơ��o�Dj+���1Z��B$��[�b?�"��'�$��>�Ym��UxӦ��gd	z	;jI�Q���J��&�UJ���H�3z�����%ꗯ�<�J���ob�Fb���sO�0Gq�H��k#B�rq�+�`��
%d�T�Jg�g'�I��"���ʀ�$���Q��⸷%I5�M�o��:q��#��u���Ƀ|��g��_O�ѵӶ��t&�3HP�!a�i������>l���ݧ�N�W�&�q)�k������ְ�W��HX��}H�@J#g����:�z��Q!��kT�S�*7%Sl&�6@����bW��8NP�뻤��b*�� ��Z������ahtjI�V�,h�B~�èbט��٭��`L*��?}�3��
(e���[�(��>v�94j!�����k�b�2��S��[+祈��Ϧc��Qm� �O�Si0�(�\hδ7������K%���-!͹&�J�~�H�u��n��?,P��j.z��G�}�����ǃ�
�y�w�G��nX4Z��l����Q��a�"y��Z��o��D ��5��}(��w��ފpa��n�Y�A"SL�h���8�Paս}����v5��e����
�G��WC���K�=oye e(F��^y<�IqěѪSE�Q��c;'�\0vӰ�$���4����H�	O����=�d��>-� J�)��`"J�k�8O�W�.O��kD]f.�".��*UF�� N ���	B�]�Yq"M���ȫ�{�l�4� vQ��Ё{[��ܫ�ۮ��>����Z12��|fw�rQ��2��*Q��B�����h��۹�|�D��~~+�p��D(���
�$�g������.�%p
W0��G���LQ�5?]3�4&U������w��Y�'u��{T�@z,z)F�YՋ�#֛<S��ǽ���b�p�`��1���Փ��}ٲ����&gܺ1HM_�}C�ˏ�8X��~��Ηs�l~s���H����p�s3�;G�J���јx �p�~�ф�$�Ӆ>�Q�&�� �r\'��6�A�'�.��re�-���`h�����$/7U��_�jLJZ-�x��2�tp��P��V�zJ}���MC�D����9����{��O %rK%R��*tA��eM����L�p6 r7u�9j�|s0bQ��`h�l^����0�(A�>T&e=���܌�X�҄UH�88����� ���L+��,��G�d��n����#��X!����E�o?,�o�R��+�����A}�ʝ����<�Z*$"b���qM��I�pf{���`�<)��V�B� �*�W�UO���fZ筿 g�LP�T�G�}�����#�A�833�����Q���.�)�*1��ˑ��N|"���鿇{��yc�^7�7j#5��*��[C���H)�V�Z�r�xOɻu�3���҆wNː�c�U��Us���`zxVE�8�X�)�|�a�X��L.�]��&�=%v���.7�iT�]�M��^f�-g���NQ�ڸ�IbHoC÷�Մ�?F�bh�c�ӂ�Ƀ:�ۄi}ݸǝ�x��ɉYo
)��:����������0u��gx1"Y��0��~LO�#����՞�M����BM����6f8_�;#��"��sÜK)ɭ���y5�P��=�i/��3�O%�}�ӀZ{H�ؽUe��W�l����1���̃p5�C�s�a[g�~�;�9�b/VM�q�<<�3t�E.A�B�Z�d	�'|8Ŧ!嗍�5Q$����x�v7<���t��&��D���IX>c��aR��"�O��^r#�@�n��)��T�/l�6��ޘ���h�x�߱��O�}w�E���#��HRѥȁ�!َ�́|����5�"���Z�,�#$�{�N-���d�?*	)�?�k�==R����
���x�0m�b��͢��FH�����t�#��/�k�O�.�3��9��*N�E03�!|#!1�����j/4�T�.LK��w����ْ�
���PE�ó�@#��)�x�_�
iJ�#R��)�f}���[_�H�e��h�9�.y��ϖX~:k����x�@;���Q�=})�|9 {,�:�>��FS���3; )��k�Ƃ�:��&Q��dEA�!�aj�k��b���C�ʞ��֢Q��T�we(��A`ldp[s�4�����R���D�34T����G�FR�V�ًZQ,;?!֮��˅���]�Ɲq�������V�H#d� h�M$��J �#M{�s�=�$C[��4څ�@0	Ps��kk)��-ȕ���Ph`Y/�"�1��/���4&͏�>fm�o��!XH;5~U�����{��C��z���W2"@�Ǻ��{�b��;ґN/s^i�a��/�GA�yH�����^d���>y��z���9��]�Ą��V#�V�P�ϵ��K��N�!�%�>�`7OKxƪ�dm�"�w�ӡF�5�l�f#D��}!�e�Č^���Q�;6&�`A�W�fZ�hs�����n���j�3DP�d�Ug^s�����FEX��+�%$q 0qBt�3�@m�'��OX����{���]S��6����;���0�� ��D4yGMn�e��d��r�P`4.��'h���]b��e%}?�!#]��R��Y�9@RQ2���|t(GΚ
c��Ir��B�]�����I��S�-X��^Y
���C,uӳ��>`��޲U�_/�GRS����6�si	s�W��5��Y	����:}z
�U���n�?Ƃ�7�;\)�.m��s�,�-a�&P���b��Zm?`�y^hn� `�$��ξ ũz���5�9+��!�����w�D��4���E���;.�s���u`܋D�E���ԑ�v)�|��w�^�������Ȣ����Ă���g|CT �����أ��U����$����H�!�-�?h�ntr� ]��K���0�-b��%��m��ơA�{��5���)v�6˶.���ۧ�`5����+(QY �KF�c����m�!;F:�:	Kl��\�?6p�g�7�Q��]�]G��Z�l����"T�k��=i���% �/�[�]���_։
M�%�Kȓߐ����fp"N�I��82�=��+Iy,x<��r�y��.2z8����Z�u;�������"so�S�����.��7/�(�2hLe,K�X��6>퐒{�-���S���rv�ƥ�8�j|�m䜮K������(	S�rɶh�~�Sj�{%�qxf���A����B��]�R��i@.�&��G�|��-`�֥�uY�I��<�|���h�x|�TO`l��5�Ԡ�J}�{oPw>M��ᵽ�p9��ܖ:��
)�6�oӵ���F6��qae2��M��a�9�L��"�{�e��� ���T�7��xD��l�����ݬ�L4oEcV75��>q�)a�?���U���1�n�m3��}�s��l�<�����K�=\1��Yq�؃���N�Ǫ=�DXH�+q[�t�8;q�'��Q�������/�7���.}���
a7�B9�cd�>���&"r��2�s�v�B#l 
Nc*��+����+=.�;hV��`�`��2������
������yV���1J���>�I�ڣ����Ѯ/��&�"^'ͣ�'ʬ3$s����\�v�dJ�>��A�#{���fsysF��=�Um=��yE�	�IT)[/���?s��/JJ��߰ǈ�k?A�聃nUS8���.����l۵�׈�-a���Ω�q�X�����'`U�/PC^�ܐ{�SY�jȔ8s�l�U7���ڿ���U��X(t]X��w�\�5�����m�|q�U�o�3^͌m�'22�7��A�_:��5�	xf���_�E����`̛�5��2�M��,���P�ol�hF'c�`1k9X|���]���C/���*)/{�ݜ�����ɵx�5_)	3v���f~a����Kv�1�B̹A�fM�)��I�v����<T�ëX@k�{
$�Fś*|�u]_�y��j�H��H#S��ƻ�T���f{U��M�ہ�0�i����Л�(_����J���6[s�\�����r�H(�7%�d�l�����}z�ʉ3;>����x�����3n�l�+��yZp����WaI�瓶/I��C�'����F>Z/.�3��>���łsB̋.2S���B�]2�������{C����F��|�+����l�h�wZ�F�������W�_�V�Q�2l����m�����*�eacv��!���F)��u�S8JL�x�]���{t�`�����`�s`�F�q���g�MӍAK?U�����ȳ�|{��y�!B�:�r
�٭�ޝ�X��c�Ml�'�yc�ĕ��?_dԵ�"��u��� ���P��rFeY���_�(�_�m�z��ʙ g71u������"_=SMm$�{���VԦd}T���wX�sL�o�w��T�#�8R��q��ɜ���0�W=Щ'��51�h�:l£���ު�S��P�0�؆i�>LfeJ�����p[9iCg��v�(����`�`��܅�2E���,��^V�Z��5�D����l9�/y�k	M��3�&5�mDFd%�'�K�L!F��Pp(;�a+\"X��;�b^M`�a���k��.����������%M3���D2���%������.K��/c��h2dT_^�C��&���{K8T�ɛ$�3�Bi����lPMv\W���XN�`{�5x����^���a "�oZ軔��.�����"���8w��Se��GO ��X��,�)F"d�{#h�w5h��]^���Kh�y1_J"��y�6:��0�J���K��S�(�L��U�F8��Yyz��Х.B�a��q8_�*��AM=���pME�E������wP���@��!��;���N}ej���O.�v%�n�B�/�a*��y;�/���UP�A 'Xƌ�ѽ�،L���}i#5 򴆿h��EQ�mKm�R`E���\V���D%1tW���H�ig���ұ����� �b�M�A[���ݯF�q7������&�nB�e��*`�M`lY���گ��lB���Y�q�eɀ,.4  F��G� �s�}鹿�2��4A�x9s
�B���T��.����Q�e��eň�=k���&!^�:e���2�D�5]�8�q0�T�Ɲأ [�v�;�քi��IRp�y5d1�w5�k����T���-?p�9+���*y�/�Ο. �nZ�Py?����!ޗ 7�����9��F��~�����|������ɍ;$QJ��d"���8�������f�ܣ4$���:���8��qxPC����q����,R`��3���mc�J;���,��3�yMY����Dێ�P�Է����S$}�֚�)9�x�u=ob�7��q��V��ĬEԇF��_������(t�c��
�aO��2	�f�s�rX6KN����6.��jQ�����
BT�";Er�U#�zY�y��#1�����ߞU�r�C�/�Z��'QM{�f描��)��U�kk-�I�i	i�{92ٗ�6����(޼xK���UD1�CO-:_�ƠrңQ�
8/�v�f}�r�R���F���c�1|Ŕ�Ӧnk�cP��I�@z<�&��7[�m����<�U�61]+�Y�Ǯr��Z�f����>����^�N4c�i�yu[��q���1Hk좶D�����uf�ow!���������L��p���ݱ�]��7Ǥ�5�
����C(�%yckt_&��~�C�M�VNU�H2f,Wf�cG��C��I�C���k�f������
��NJo*�s���˝���i���tKl�������s����C�<�N��`1T�Vz+"������WD�N�ɞ�QB�����x{���.y:V	������u�L��>���I��3�i	�<�@2NA��#�G�޼���>�)�>�R�͸�}�D����ݩ���y��F��=輽K6�{�G<����4a
��y2b$ �Ck�q �����eNЂ���{��9,q��F�p+��y��QУ� �� ���)F�^�1��΄i
=��&�N����g+�6G/_k��X73�~-WH��\<����P��m�4o�,F�'��<�������:1��֏2��əi�Z:�?N�G��N�?��^2#�˽g� �$UR�+�Y�kiݷL���ϸɏ�:��[!�.Sr�Uu���u�`�`�tSF��D�wl��HXM=��9�C�	���Y�����C���4�a��wj�����9e�߲��	1奬�@;�ʺmw͚�k�/���-�|Ɉ������ b���X���_�>G�.�%2P����@��F�[���"�Kyg�٠g���v�6`h.���������[���� -Y��(m<����[v���t3����%#��m%����K&���e�iz�1*�kw���"M(�����!�����g�����Z} ��A�r�/V}� [9 c�I�e�-^ol����pW��)K����߮wT�H�;6o� ؟�9K28��ɘQ�q�b�Q咽	�g����zl�:G'z��Յe��h%�@��e5�����&Ig�������o��ףcI*�[7���q����$�G|�@˪�f���� ���C��qU�n������שO�i��=�O��������le��Ka�w\FH�:c�|���(�?�D�lXVC��G.���'��?R<g��D���s����g-/����A�Y��Ɩ��_�'B�]W�����SȻ+��t�?-�g�d���m�������q^�Ĩ'��&��qo������P��c�!�o�I@��9��Q��^=`�N`��ɫ�������e�(������շ'���%A�bdx*QF���n1����eF)dt\�F�X|'u�1�ʔMK�8Vd���'s%�ե���ŘFB҃&�ED� 2��խ����,Zr�B~�ŀj�U�lV��l��jmi�K#���k��S��x �GY h�	a,e[Rk����WJ��atj���C�r��A4�xF^�I���Q� Z؅=�	�t��f�+R��9����m����L�=���]-��0����!�Y{j�z�m㻰G'kA���/ܜe��.��q5}��nt^���/ӊn%����7�� [$[E��!����1^Ew6�eլM;�d�b+MrW0���@3�m)�=��&3%o�'����K�#�	�EM+�k��+U�vx��'��e��]$�_س�`����k�=8Z���R�c�H��́5Kv�<��K<!��Z�%�ldX��_3����+S���sK�rNIFTz�d��
3�Y���@�����������:�8�eƀ�+�L�F��0ku��j��ֻ�\�n8B㠚H�<������j���W[��km\�5���c������i�!����(�,'~�ރ����N�\;�A:~H�ëF��T������Yz1=�1��ƫ��T�p�WCF�R���RQ���!/Za�A�]��c�ߒ�����&�Ѫ?����\FP�V���Oѝ�%e��dr�"��L#O�5q"��U��!�е5�{}0�`B��@Xr:}��.�RSU9�\�C�X)�8�4}'�+?2�KV���na5��l^Y�6�E��2y�����6m�EY
����3��׏s����d%+����G�������Wq(��Zî�E�%G���=�1�|Zd���a|�z�Kv��J������/V�n�ܸ�k�����'tx/��nWb/-Ƽ���u#m�IEU�~�֕R���ہ�9���.;=!��*�7���ۆɮ&"��R�������bkqF�hF*b�-���)��g\K'���%�6��I�ƈ�z��=Ջ�w��@���ö�0<���vr}mJo`�y 2�ڤ��=��)�˜��o���2�d�흪=.�P�P�QվvAQ���[~~1���~f��5/�ַ3��_�F���&R:���XZJ��7�*pp�S!��捄ł�O�P��:II~�v�+(�5 U��4��7֣j�����4���� ���b0����7�3\/�F�;-��
��4эoǸ�L�zv� ��Y�/H�)�m���Y�!�~̛ӡZ�ܘ5�j���Gc����.)��oPH̞>v�_�{�U�eWGZ�./K뉋*�O��3��H���*!٦#��D��]K�'k���g~:��LZ���i7'<��%�1��ƍ�BN��L��d�C۪�]�S�I�ga�Re���lwl��0QfX�&�ۆ�U�Q���֞@��͎���c4*���g�-MCj�B���g�[��kL��3��g�J�gk;7�lF4��3q�u��o�8�͎�i�v��'9 TG$o ë���Es5yZH"1T�����f��C2�<�{��T��t_7�,]G���=��2~cN>-SLїX�U}>^G깴y��2��XE����J���b��Z�z��9w��v�8�Cz����8XsՐd6��+�.}J~���m��)Sg�ʏ�d���Ò�N���lD�� �Le� .����{Ł����d��붒93�Gm���~��3����{�tGόf�"����]�q���C��ٲ��m��H?��ȑI8%�ɁG����a��T����֡}�Pk��l��CB��T��K�Oc���o*���"N7�{�odf�u�d��;�����÷h(Ś��QC�>�q���zB��m��=CN���_%[F��5�VLJ�4���,}L��0峨΃p����o�.����ϛ�C��`ȹ 8<����o1�d���-��D�k��п�X��z� �D��mϘ���%`Y��Ҿ�;����	�f��V����Y8?�?�q!�}ؐw�n�����(S����D8
������~�dѠ�p�2J�Y�x���}�_V����0���;.�x�p�?ĬNB�� �灻U�S��MO���TVa�Z�0z	��+ZkH��M��_���ý	7
cX����q�mF���m׃�྘�?R�7r��,�ñ�/lT����ؕ�!?�0�Y�D�);���7$ա�6#�]f��9��lF�2��D3�9#���<8	6uډ�4A�{oLcܾt�`�R����1@�z"�w5�z�B3��?0&G2������З�e��M�Ʋ���ïT�bC*y�?3�:�O��eD�(Յ<���$�Ѡ��f��*G��:�k�n�Vt���Oɝ�����ƥ�x��ϒ�Jnw�9y$�*����]Ԣ����x��[��!���^<
T&ݬA�_G��]C��K�@���"M���u ����ۊ��?u`���4�>�C�j��B�6��K	��W��/�'/�؉/톴� F�{A����o�葮�4���$ � �pyAw��V��ȯ�o�Ɂ���ᬯJ�o�y[���(g{�S��b�ҙg��Y8���8X�+]�����TZC�a���ͷQ,�`X�
!�\�(�)���7~U]w=��w���.{� 9��Ef�j���Bxi�Z�V����� �CM���n���2fx�f
�As�O�t^��o�R$��H)��l��^� �v�0�]O�î{��q_�������M��-e���;{1c��;���;���L+�jL�՜�z�/�24��u��O�]u.i� <9l=�'��M�����Y)z4g��irrL����+3$/癈�e�~��3:���~�'��pbxo�w���Q7��E�z�aR�h��\��`7�!�%���<+gc]I��	���&�T�o�3�]�l��L:�^�Y����<?���hޤ�qe�6���P^���w���,*���!ɄrkxO�I��w���*�yw��t��9(���l��i�HQM�sc*n7k嚭0R����H ��a�k�u���#A ܤ��]3�9��ma�_s�V�&3AɚkP$���J�K�%ή����P�4���Pp��ARK�<�>d����*�	����J9��a�1��R2�#���"�V�`�* ���Us�rx�� JN�]|�o�z�M�&M@�;� ѩ�e�W%��մ�N�4�I��Dt��nuf�s���Y�����w�xF�f���ׯ�(Z�c�I]iqs�ޟS�����&�$}�Ä|��] �F�
�>"QP�?����G���=�ʒ�� ��|w�(�h'��nϮ�}�P	�2'=p8�6Ϣ�%L_��|~��_�$��~H���^ި ��Hm	�`M�<F�$��t���@ղ]�t )u�>R.�o��`r��g�&e�OO�k�����S��4�Ix6_[E�W�eC�k�ޠ�wOl6T��c�s?s(�<�zu����р>EٗQ"�+���jC�&H����ޛK�L�uY�Y�R��3�`Nw-!�}������U,R�EPH՗���s�Q;��:��<�1�#E��Y��LS�	��
�g�A|m��g��p�4\2������@�>���f�����N����J-��9�aaG��OoVT{��p���62-=�|�4V2�Y�%*y�6l�Ә���k��r�Y���IMcY��r���U��\���n�:J�܎e	Z*�3WV1�hb�+lDE�����X���կ�5�)��^�{B��N�8���y�-*��\��́6� �D�7�~�׬�	c�����h�<6w��wT: �j��	@Y��	AsT�;���;@���!􆌾�޸j�b�ÁJ? �l�qj�6eir���x�0/+�J.�IoM��8S��>
�E����s|m(�t�L�W��ʮ��A���[�A(�ɞJA�Z��e�F�ϙٛ����Z����	Y&�"�]�h���3aH_BCH�#����I�X�G���N)	zI�a8�M(!a�7�������;��������4��+;��ң�
��o]G�1b����˰%k��\1J�X��H�N�,+O� �m� Ҽ5�)����k���F�^ y�UrNq놐�+*8�5�2������jS�e�5徎C����X�Q�0a��>���j�z�j�.E�-����srzP���ǻl׉��dEkn�gЉ�7zb���hW(RE��J2n'����`zُ&Hl�*�V�G�yh�A��ٝ�D�?*�th���3pö3�pBn�D����A�z�؍:!�E����V�nu���Q������(/h_q�UJ&��/qjH֌���D�|�=��F�����(�Z:eW'5m�q��ȹ �6��\C�TWa��<(w����Ye��2���;�3��u3&�C�K�nr`?JC�K�Nv+��OL$t�@��)�z�t������̐z1�N|~PJ���L�W�. �S~;��3_�O��?�0�w�X�@�������YrTk�>�.L#��"lN������#�ϖ�C̭\+{0m�!S+=���
���Ȉ#Iq �zֵt��e'0R)�fF=1w���48���a�x�\*U���1"��'�-j��!���u:�}�Ά�z���KR%i �R��ݺU����}wќ�q��ds��ο�W�\o;r��)䮛r�6���A��Z�0u����3�<5��p�N�Ő�����C1!��$�/R@3����$Kn�P7]���d�zx2rU�w��5��؅w;u�<�vj}�7���8=|s-B��I`�v��4�@��V�B,�R��klû��,�Lz�w�qt� ��C	���U��7iMb{1�:
V��l���� ��V�Oq*Wl|bӖ��'��:�qZx�u�w�<�Q�����m���"ޒ�� a|z:I�����#)'����$�T����z%}q!�[�}9�%�ǣ=i)RI�t����w@e��GZ��4���G��?�]��^$�eL0Ht:Sk������G�=���n�Q)8�'���Q~�2\�?@���ܙc�@%{�׬%˾�4�uHb����
�/��=G*A��iħp�2�7w��[P�\�܊���(�XJh'����F��+@z����[V��O����#�?n��\d3�D���>�	�M��pr�i�{���H��E%��F;R��/^���;:I�押mS	��to.cի(�攸���b��sј�����nr�>j�v�Lj���pr�s�HU�=d`~��D�,�^����\��V��y> �h����7%o�}#:+E���Gk�s(T!t�k��,�+��ao��-x,	�&H�(fS�����]��6A�ue��"�B�1��pڻ�����mumgOi�gJ����F�5$�Ϩj��X#=s�M!�	�<�4�J�����I���z3����A��ɠp)�3��ݶ��L�Y�	��?ʤp>�&.A�6:y��(�������h��xE"S9�!mS��Tx�9n�r3����E�zQ�+\7}N�x��:�­`�KO��eF���g�ּ�_�]�E�t���67Q��-^��&���7�ۉ���e���n�wV��x��GY�F�b�*�����V*e�s�d�u�mY9q�A�Ӿ)^.c�ԱZ=Gb|�&\5�7ݫ9�F��E*P�<9��"E���禹/V��N�7>͌O��(<c��O���d'��]���\���c��2Gǳ��I$ֺ��[o5Lt/�JLK�l`2��;� �f���,�'yc,}��������5���ٽ!ϥ@ɻbT����#m瞏��d��UM�rb��fy��_��g�xkܠ@&Ă�1�^=��,�� ���f�e�QX�W�i�W��S�c��ä����0��,����*@VT;��a�(i&<N�"n��&�R�a�
���=��(�5K"i��$>���\q @�A���5�2�8��O�p���Ɣ�=`��.'F��@U]��"T~|.�ԯ2T���$}�h�[{���Eh�H8� @|�yu��y_�[/�{��%P�Qdt�ҵ�Zv+uuQ2��3�ҡ^��%\<���{���	ά���(�J�ׯ�xM]	���]�:6?���v/^�R�Y1�qH����?�O�ӁՑ~���:�"P^$H2���{�>������Z�W!/��u܃=T��k3^��`u��b{2���h��; 1��2ӎ�+eT8[��)O�p���[t���'���ĜF,^���/\��Lx
�8h��47��ѿ�F���4��Z�I���˕��ьd�]���˂��M��S�'w��vA�3�6�HAr"CL�p�w���P�n5r[/9�`R�v�H��ž�
��A_�ƴq������FPG#,�R��`�]x��E	��9��~�6�����yi<�ʺY�vN������C���n(4�O��놔z�<�F"������֡���?rv�?�4I٫�N[嚱���I!A��S���H*�^lk�0�,c��I�(���iq�v�����v}������d��
� #V���P����18�`�=;������ҽ��� �X�ں�zKcdeg.F �����fhGR�nk�fO�!��L����62��E�n�!���qpU�5E�|̀!�^��ǫQ��)ٶ�Ka��6�
\}���':K�l�(e�z|�I5��u�7.�:PpX�τ_ɸؠBq��'���ZԚ�������aAo��)G�贃{}kpU�lȔI
��qПX�089V��4 X��p�:�ua	G���d�S�G�cs�,����ı6���<���-������^��
��qA3�eYbv��N'l�cV�K5�#2j2���V=i�*�C�ɗ�̝�����A�-������ݬ�����#'K_�m���	.Kv]ܨe�Hk�:X7��d֧>�+��� �Ÿ�P~��ӑW,��<�rɤ"�u�d�Ȉ�8|M���f2��GC~[M�t�w:T-�x�E@;h�~�:�H�]"K��;��)���/?q ؋~�$��9Q_��2O��T��>�?�����v��B���X\�����������B���wu.��:��NKD�:\<8�$���==/)���+߈I� ě@�<ϩ�F�I�>�m�~����KL׀��ƛ�Q���sѐX�t����9�)�n�tԽ���E�P�e�=�o���K�7%.*?L��h`+�{a<�`ž}á}綠�y,��1�{L��8��p4~)\h>t����/ڠt�3Q��������gK��7)@��z�)�XB.'@\si���o�>4UA�<�a���+z$C0���9,�b�CǹeG,���6f�S	�P�!ӥ����we��M��e(�w�x���Wؒd��h�_� 	i��ǯ�4�&H�S�DR�~)�0��-	0F�%P���Xm67H@�28chqV�	:$��E%�2پSgi#DB��3  ��w�x}0�������}�p�+ڭ1��s`�\����C��k������9B1-�m~��pڏV�J?/b�MX&�%<�m�Pw0��?Sъ��4��)��t���`��T����� z�5:R[	�r8�;����J�:k�R�r��~�ռKH���SE�X �N1sO��":�:ҽ��Sl����X̳P;�.Ke�?M$֡-�f��o����`�У��1�C	*:f�u�6~���1�r�/��R��7���"!���jP3imX0��Є {��1YM�E�0K�TZ48a���E��z#x����»�.�:A�UC�
Lq`ƄG�$�^~�)T����d�� ��! ��L^;-q��e��P�*�I^�=Z`��\Z{�� _��g�=����@{^�0t�x��s.ђ�4{���:]�TE��4T+���Û9 �������תc���:� C�za���I�/ 1���NH�tTX�9���u��\����Dv�ӆ[�(��" �#p���Ʉ���ǂX�f�ـ{���p�Y��"8�Ov�1q���9_jG9�lQR�5c�=�^��B��(l�|DUJ�������tGy��/et=3;c�_2{���J�/�[Q�3;�g%��w��.�z���z�����e�qσ��'�>u�S��Gc��V�s�@;˥`�	kWt�;?�;�ت^Q�/�}�,��K��)Ԇ����0r��:���0 ����s�H���X� 
�##��ýx�N���`��b���2̗s�!�M/��|�V%���-��g��l�_�s�w�ZZ7J�`���M�ߖxeE=��0N��,��`],ק�1G��,��Y����\#����d��a��(�����t۫���Zq_��t�"iuy�895��c_]�}���xIn�맿��6�&J�L)�*zl�� ���p\��NxM�=��6HJT������5����}N<��h����-i
������̒��l���̢	�-�F���q�]��T���;G�Ok��&9�%b��t��Oh�
H�� ��wghő2��v5, S������#*�ߛ R���'ek% �r���q*��.P�91B�s!jF��?d�F�ђ��Y�����-
�6ђ�`��:����cE.�����YU��`�Xu�M��i�򦝟+I��b�I���Ș"\+�<���ӱcS�_NB�Y5�{s����J�HUq-����J�2j��X��t�)���AC��n8�6W,ws Xw)��o�h��t���'�F�>��������(�F��MD�#�˙��os.\=�9�,;Z�T�T(&1�J���W#Xm".xSTI�k�$̃��>Ǻ���{I��W_}����A��M�Zi���Ӹdl-��ͳ�r~�>�;Zq�Y�hN�`�*��� ��+6�"�gjs"��N����MЮ{�ۛTu�����@�{����L��˖2:g:�GԟD�%�;�K��}�ݮ��%�rO�ԟb�P\���oxo��ԅ_������YW--�?� g)����-�  ��hi;����Z�NO�';Ϟb����Jfp�DN�O&E)��8���a=%׹Iu_wY���]YD7��*�"��9���G�x�G-�>>���l���vd���kj�ҋ�@Y�����Џ��Üw/�D,�tw�U���_�q�-��]���~�Һy���'�� )�^������ZİW�����P��!צ�"���eA����7�Ո�^K�[Q���ᖳ��-,���<L�8���5J�@���$�kV\�8��z�e�ӫ�eH:M˫;i<Ӌ&σR9�b�HA�R}�n��`C�X��b�4C���B��RjPV�ׇ���L�6�cZ��f���T��S�3�	�+������pˏ��P����m���B_�74�Lg<z#Y�A+d�MK)q����S���e�@}������(#1&}/X��@vL��
U/��������tt�9���[BY�۝l }��z�#��0��.���+^�Q��*�L���Z�:'v�ʘA���˃~3�Q]�R�����M��N�I�eu��]���x9���k>��i
��7����l�j��04���`w��nvR�Τ�u�Hjzfdf���ޕ�B>�$Τ�"t@����Z�>��&�ϸZ���­,�<ֻ�L"������<�)e!�|�L&��u*Y��$�2P�;�u�A�Q������i��΂=Mw���&[|�%;]���s�+��#w�6�<�_1�Ǉ�������vt<H���WN>RR��+�f�q"�*ۜν�XQ՛=�qs�6\�1P�?	ux��,���$���=_͏e6s8")�V��7$���N����U,�>ˊm�F�����Ayp)4x��p��E�^Up׉�5�S:��w�B ��-�q2yUh}�� @�G������DZ��	Q<A�b�V��׺�ˠ"�y�}7]}  �o�٠�K�V&�n.������j�z����`�d��i8l2�*r�N�a7b�qoNvW��z����\b������ip��ǉz����I]~8�1]��ً��m �n������F��A��� `9�!�:O�rÁ�*U(�LҴ� *�/�@��'�)�>D�hY��^Dӗ��}�����_J�ΣN�������H���ߙ��6<�syߞ!�;��*b�U�-�:Ǘ�_��mk����'�
�	RV�e^���v#:�XeS��Zggzx)���ЃM�,<�:��|�׈��n�IZ�3P�J�T�5sl=�.����G���.3B	�:EZIFϪ�}=](�,�t�Bj\ZcJL���6��@|�=�5�
�����������;L��Z��PB�Yöm	D���&y��
LgW��N������k�W�+�.iw͕X?�hK��?�#�ѭ��h�tpz�A��޺ё���D�
�(�<A/�8�+F��9�*��Q"�@�^�i�|VY��"~_ZQ?B���3��ϳ�?.y�Vk������?�U�C����c��c��d���1K%X��ۢ��h����)q�7\�$�?��|av]���M�@#Sx�I2~fXnޤ����F�6���9�l6Yz2(���Ôq��k7���͏��\�I�f�"��9#9;�_�M�\r��"T JV�"��eS%z*b�����(W���K����A�[�)�����E
)]������D�����+�� �e.h� Ta�!��j�E7�;��D�
��D��#k��g(h���.�<q�][�ݕ���6z��*���y���ʨ�I��� ?�
g3]lvU�Y���/��g!Ő҈�ʤ@5� ,�VCę	���-�8���.^�	/�DRA��I�W�c�5���b�5��"� E;�G��YO�〒�@�~�U�d�`-e���� ҉�:�XO��[3�X��T��� }d�G�����j$�k��.K>O3�����A{��L�mӡJg��oori@���䙦9���̝|1�(Z^q�Ę�������M�1��VGF��U7dk�+�u�T�lPGc]��xbc�J_�J�?�v.\����fכ�c�E/w��Arw�@V�@]/�3<�[����|� 'U�0C��T(gq�z�K����s~�)�	@�5.h�9�2;wn�F�:iRi5P�84)�~���m�7�2�f5$p���B�Fk�&x�� qZ͌b��<&}qmE8��-����_�R��ѫ��Ga�|� IYX	Ms{�#�9�.���:Ws�*��U%���h��+��^�2�]��'	�c�"�O��N�O{;0ʒ/�
��\ ����&�
Ϭ��AR]Ө�����2֚����~���9p������h6�.��P[V���ö?����M6��1��{�*V/��.��Nn'Pf�hU�"��f�Y��4��
yJo�N�5���L�Z]	�K��������8W@NO&�k<;�غ{������t�Dꃕm��*�*�;�a-5C!��v
��i�z�E�W�sv���n���xLNH<lv��ȿ�b:�<�g�:�, :�jfy��ݭ:x�7\Ti�7���NY�Si��tNM�-!��w�ǌt�(=���:C
�
aս�(��1�z���B��Ϫc��T�����G*`��pI*{
�G�8%�+=t48"�� ���X�'�a:�l�A�?^��͐<��s�ZPP:��T��|�c1OJx��#�Q�ؖP�3GMI�k���	QN��=���l�
>:k�����ѻssn�~�x��c��Ⲹ|5Hj�<X���',��1T
��r=���Gb�����7�m�� n��.w�]����!�6
��~��nr/SV%
5��N��� ���`�=дB���C�<�b�<��nY�-�/Y���Rb��Wϕ4��:F����f�JmF���/�v�\�qcg0�/�(|�
K��ɈH;V5��,��H�zAm_^��C��;q�im=h,}�sn2������X2�W���F2�����3�8{_P տ��6al��J�Ѩ��9�m�����\�r�|;�:���'\�\2�N	 ���[�vL��<�$�#��A���J��Π�U���� }�:�Xɼ��W��%��O��1@��uHY{������G�C#E�v�C�w��:?�4�\��),YgL���@��O0���T�YշU��'�v`8)�mW�L�� �!�s�
۪�E2enjh�O=�K���M�J����9�	3hb粢�aks7��š����wg�,<A	�g�TP�FW^J �&��~��]I�|�M��B	Ȕj�(�OX�� ��q �<Z9�f�� �u�e�\��.����l�ӧ�by��<���J�dc"�!l� �� x)�A����~c�Z�s��R^4E^�!��]y������m����zt�E+U����;�K`kKt�f�Gv��KR��@�G��6��ʗ���\:��3,$��*���yg?�y�SG+�7�a*��S��p��������Z��ÕڸA@�H���N"P$p`�D/=���dI�JVaڨ�c
o�h�8�:�-Y���?Ya5���A��h��~�ֺ_hRyw�F2���!l^~镦���6�7SP5.x��8�
���&{���]�ǒV�ŧN�L�2d%�4������/O]�v���o�,r��A0���3���S��*\d����Y�rߥk쾾l$z��fV�I^���s`���9��b���Ǘ��äH��.�k�3韀�-6�g��	�b\��B2�P�e]����v?ɭ2����z�~=W�M���}v'�'��4��� �� �-Oy��������9���p�}��tK)�S�� ����nF�U�=�F.���!��>���&J�C�]&M� @,�>R־0AH��1�i��Y��aW�R&���f)�O[��@������(���$�aӤ�6]{|���	��4�7�ű�����~;-���D)����>��{��t��C 	�ۼ3���SgX	B�M"�S��q;#�h9�բ�̓���o Zד3 $��	�|�~�ǘ�_4�v�~����U��>^������3�qL`���.�#�h8�>-&+��S� _����Y �7�K�ӔO��ъ/@��B��[��:��U���G�{���7D)���34��NQ؀�B��֗�;I�����P�7��5���d�#:�/:����W>����8�]����G��Jz��\��������_�JSj4�(ob�TD����w;+Q�q6e0w1<��
�Mf�� !�9��m��5�:i�U�:z�A�����FB�S���쐩�G�������
Ώ� Aop�Hu'�R�YY�iᲃ5G���E9�������)�l[�P)Ь�o89�+�W���I'oV#Ѭӵ�	�'񨂑��7�?�:����ڮp�H�� �c��?Ɵ$�!I�3���u�,h�rޞ#gr�:�?w����n���g�� 
��Z�V:��1�ZA)�D�Gk<�>�-��H�.ao���@��(e�#�x΄|�Z�H����z�P�6�aNY�����xv��~J������
�V��ڨ	��-�1��~��U��(��Ff5zfe4U��#�p8�P>s�at��J�l��ƚI��!��i�"	ܧ�o�}�gLYh������I+x���_����=����ӷŽ%Z��lC�lN9���RU���{��kY1m�F�S��M�d��3��|W�p<��wׅ���;$�K����]�U?�K���$O�SP0݉j��G����H֢Bۗ��z�\i;��d
��y0��I���o�`�OR� A��GNO�e7t��`N?�ul6�<��rsl!dֿ�x_>�M��G���B;����S�I��
����V�v>��ß�Ē\�=Wǹ�\�hS��	�1����ér(Yz�R0{�(���N�g��O*��pz����L{�=�@�Z/Q$��xM}�).���c8��g��4n����j�c�����w�c��֖ܘ���t��J	��
jЌ�^��^\m,�z�O4[6Kg���43+�0���U����j���%6���镫�R�K�wu��in�)�N�Su��X�Jqn$J�Ԯw�$P.+���XD�T��U����1JO)n*Ju�E���`�6� KMc2��Y�������AJ���:_���Az-	
�p����� k�\[�\I=/0�V�}ԐO�Rx��'OǱ��d��0�_w���{�����=�S��QdQI��n6�1���VM�<w5�.N�ck[���-��������U����)sx�Lf��y�~C�KŚK/�Ω~�tX�a�	T@`����$4�8԰]��p~>T���s_k�o������I9��3�~�`�7�XF��X��8%>pFR{�Y�[_�Wlt e���<������_�Q�.e:��W[����4�Wh�_�C0�kZ3��)$�x?��x�;�o�נ}�����S��ߢ�����Ih"�P�'��u�)�Cй����6���^#v%Lן�Y3	�D��qݼF�qmv��/�KXy�{���l��c�o���h���k��w4v�`�>^\.��&�zDZY�b)]��j���3R[�b��J�['aI�$����O;�.ҫe� ��K�O�uj�_,c�
���X�=/0v?�B��>g7ȡ��.���4��W��i������x�6D�K�x�zם̔��,���%��⸟������m����>f���Dl+��������B{�lW� �2�*�.'���p�o�����i�N���A�C���g��(�κ���w΋���;QR�:�EK�ݑ�NB����o��ƙ��O�Y*w�)�ƿ��c��z�B	1��N3ْw��[���~𠋼9�������v�#Y��t�xs��ڎ����t����GO-���&����t�%
eUەZ7Y���TT���6x7޷��~f�DS%�G������	����-]ڑ,�[9	vS�Yqm�"4�a?=C���@!�1��������^o��{'��ME�?�*=UA��9����*�O�P����Ղ��J%��M3�+ ���]f�~�� ]�T"	8���ߔ(�2,A�������kmƪ�C?'N���Qm
NJ�ٕ�BEo�}q��mҜI>�Łi3����S�«N�+7Ǖ���혘����|�ͫ��G��3����b-c�nd?DռZ���Hx��u>C'Rdq۴�����7�K�Y�@E�	��{G��{?aD�� ���6�8�����2�;�L�rWղP�1���m�)�F_���"�O�1<�8���ҳeG@�'��ܪ/�b�o�=ɵ�%��)M�h�3I����D�4�J�0c�fe��8Bkέ�1<��F�l%^[0Xx�8-�Ml��2
�D���IOh����̔��!2M`�<�L�s�������܈~v1�ڼ�	?-��=�?;�,��4����.�� ~o�a�p���\�d�z�k��ͦʥ�;2Dޱ.�JD����Mˎ�\x�B~M�p�]�tl`Ι�x� ��.��V�-�,�
�v�C�@��&�F]"=���>F&�,���<]������N�D?��q�>�3�.=@��%,�2�`��u��G�������k��|���1���Z��|۞Gv6�F�vd�H(�u'����������;`��\8����樅�.A�BJ��i�n~�1�l�:$�=��6�Oz �3p�)��N��M��,I�٬�$��<$d1]�7̛�x���VY��8���sQ�؀��_ a�<��P�I9����[]Ep�[R�އ6������c;0J.\xվ��+�!���R��j`f�����N�Ϗ<��J�G��u]��3��"iӲ4��F���9��eP9�/��}��,%~���(jzӹ�o���-㫂a�ϒ��3��ȾP�d����c�Z��=V�����ԀB�:?���>(��o?�m�3��x"�9�]���>U�em"a��\V@,�ȝZ���5D
�����@�?�"l�7�<������&<
p�o��1��m��n�s9HNJ��E�M�@FaK���,����e�S*YKU�l@F95z��\��%&{6�A��6�6p��R^�}*G���6̌�lF���	�I�m�P3ѿ�`�`R��U`��͏���F�R�~�����2�^؛����u�]����$A�����ѳ��a��æ�x�����A�5�-z���Z�ol+5��'�D`Kit��w/3Mb4��" �-�o�vXFo�f��	�,���}�f+����������y�M`��Kn��Z��k�h։�MO���5��~ ��c�QЎt���֭WC��V�=�J�Ĥ�E�y�`*����;8�[`{Eڇ�a&�J0}v`w�%�RC� T<F��Ɨ�B��FO;�ss>�طhbl�,2Z��m���.�����Tx�E_��z��0&V�)z؅`0pV�ء�'��9B2~�x�QU:7�'d?���7��j��6�Ŗ�F���;��E�^K~�?�c��BU�de������2����Mm�b��<�I��5G�`����>^ޣ��� �kCU3��U�� ���Df�pJ�
�� u��ƚ�P4�@����+�&��0����S|A���9�]zEs�)Mm��Q�*�Su:ĪH>��x��iו�ܚ����X$p�������DG��,�S>{I�����,��}�0$)nԟ�r�C읽�R�5�O��9���k��_f���}E����i$J�����7���,Ʋ�g`��qQ�_�ܙ\g_��88���z�u��$�N~��i�j|���`es7k� ����V&�b��$��]�_fn������D�I�Px�O�2�1}���[zqF��,v�\?�Å�3ә���~���%���f����Sg���6`O89��y+8Gd#	���,88h�;�o����)!L�dSD��g�1�D�߁a��b����ԯ���ZE�P�yr�Y�i%Q��Mc��-Y-|�q���O�� ^���n�r*ٿ��-<u�sk�O�we��,wg
t��~N��Ix���u���Hcqmf�Ǝ
���mnt�BM��/��j=]�r��nBr�$:~X���=8��	�ld۸d��|��+��n8[p�J͐ �Vи�3ܢ�[f�6�ї:��#%��e���~$/��R+>���׹s��%M.��C�V��i�	#�k��O�M���v3�Dǧ�8�Sc�2��Z�&�T��qEu��{�)�Inlv�D����_�g��j���#о�x�ߙ��4�"�)�T�J�lc�pZÈ"K�hݭK��G� x����t�!13hb*-���$�m�:	�e�y�$ǌH������x�X*�΢b�d ����l������=����jo���j�S`	t��p��R)R ��b���g�	";�\D�>f���N��вs�Uӓ��~C����ӧs�=c�L�7��;ِx�JH��,H�b�p���]
j��\w���7�T3��,N�%%l�c��~�g�����$�EX���(4� �L�VM���Q�V�!p"��D럟[>�Z���^(?ќ:�>G�����x���z�3�S��Z�gs����F�)��l^���B�^Z�y���9'3����t��"���ڴ�����/Ͻ}�g�b.ot�9��|����wOnBt� �`���>�]��_o��痌�Eu}��y'������΋�q�]�g�E��Iq����m���O�=A���3��/�id��$~�
<j��f�6�n�!�v^���\�J �y%� Ɵ�ˤ$��� M��Y�0h' ��;�����g��������_���5&�����uBg��*$�_G�:��J��R&�ı����O W(E֬�ٝʀ���z3B=�oIꡈ�W3����ǃ�,g�ƿ���T!�ٟ�Pk`��w�}�uUK3�L���~���ěg쉣���%E�������q�uN��'GaK�뱡&�;�sw�C:.q�i�J]����$L����"�~i�}��O\h��p�`0|�E��z}��qBʸX���u;����a/��9s w�����.t���m�j�q�
�¦�wh�8���f�B-[3m�"L�M �"�X�oY��]���o+ܩ��e��q������*_��eZ�����K�9��<ю�c)j��E�-K뜹T/z��[5b�J��e��1!ʉ�"	"Ry��.��g*p�t
W,���J��;����65�/x���6���}��X���m	�2Cb���0x.U��6Y/lXi�Ъ'�{��(wh�~Q^A�+���Ň�����爣��xW.��'���n�>&����&7�%�c1k���Ŷ��4L�(�4V�U��;��S��t]�6��1g�0t2���}�J?�XV�����i�q������V�&�Ϥ��\�ϚS���2�ݥ�$��i�h.l���;\�7�H�Lv��PG���WY`�Tp`�_U}�&�����-_�eG�����.�O8
B��	"(5m�����Q�T��M���׮j�xl���	��i+��z �E�P,;�l�f{Kw�k�(�>�d�\�����i3,	��_�[U�]��g�~���$dY������{?��e3S�[(��|j�1��Җ^�kI��F��r(�^����lĺ�gU<:c�C����rMWF���*�#�L-۶���-��!["��$��F�e`v�s��F䏈&��R�?����� ���.@��[Q���$����[��Us�1�
%0$�aI^�%�Y�K`�WL��@��Ĉ����r�Նd�tE	J�DND�}�����d�S�v�Oy�[�ݟ����k���!E��g����-���HWy�v��8#!���|� *,�{�Ft�k��TmpqT4���7]��T��H�k?Z\߹M�9�㯜M^��	����X�\%;H�a�F��",/�KRK��,d �"�p魕�;�"g�ZQL&��}:Zq���d���̾��P\{ރ�{K	`Rz�a�T�P	G�g.��!�a��Hɓ��au�fF����Ên��ϡw=�����E���/@w���zc(����V��f�7��$�L� "��0iז`}���ޕ���s�XP'[kM��KKl�]GA`<n�.�: �_���-��_���]m9�}���w�?c9��g�0^��=ǒ��6c왵�f2����[�+�u7�h�j���qc�����g_��Q"���<��$�6^I2]|C�Ox7ǐ���^u/������PK�U?t��$f��)ĕ�=~(�/O�/��aW�ݴ�x> )�O<��"Z���5f=2�Z�S��Цj�=OǑXe�Q�/�|���&2��H+��g���XZ�NRl�~+3�PH�d$���:�M�����O<�ooat�ڼ�l�U2��z� �����%�y��K[\֊ޱ"5�=��(I���?��M�(\M`����/갤�JE"���vc@n��������?^�4Y�e�Lʆ��7 �s��2��i��xҞUOeQ��I�y.���:��V������2��ˬ�D.�X�~�v��_��k|���7� ��C#�Z��,�b(�,q��t�[���ڂ������wGBD��>�o?�!�;s�XS����uJ�b�45������tb�5D`�e<٩z��}%�����ܔC�PY۟��o��st��$��h�K��jL���m�Jz�a�H���1�Z���EĢ݌�xm2?��z�s��3���'V"2��s>���mmu��_~,�E���R��э�6�*d����
�ݘ�l*-h�~�ٌ�#;d����p����U�a~-�Jܞ���f����������d�h稞�d��#�@,��,��z�A�*��a)&��G���z�=Y���e
�	��!A�h�!�f��b[�D��ݏ���IVY4��П�G�$vB�����U�ք"��M�F��1H�q{��"��d�0D�t����$��rCw�O��Eo�:хQ�!�(��"f`�)��Q��!y6^f<������Uf&�+�����Oo���Ŋ�|���k�6�7'��x���^���bꚐ��w�ѹ�/+�!�\��P�`�qw~K�R��m �;W�n�P�G����Wu���<To� ?�n��;PT�K*k�|��<ӽ��x�B�]��6�>�TQAL��'oLj.k�(�h> ��Q�Ք�q���a�6�����^�esGj��7jv�r*������H��8������p�9�;�s��e!��_u"4?EG��E(�=4�����&��_A�+�K���F$��Q﫻/�Fu9V�|��u��K�R�0�u�²�E��9=3� ���$�$�9^��f��D'h�M1��6�]#�[l��7�d���a:��v�SzŹ��P�[��{F��{��QK�7^HԻ�JA��)*P!��\۳���2�H��	|+�,�N��ɼ�Y��Y��R�L���ڑ��X�d�{�������pN%��
b(i_�����dt*�27Q�z
$��B�-O7���c��(�z�u~�����%V*�
c�9p�rڳƝ�;}C� $?}߇�M�a�V�y��@/��@ ��J�(cN�(�����i�U������0���͠�#�r�/ ����G+O��$��~w�F�t!L�5�ZY�kIߨ�|��4�͞,�G�Le�N���JG0��rB���ܘ��*!s�����|6>!ȅ�L�6z��,y��~��B�8���s`pf�:|��:[�W���G���=��gq2x���3�^�e9����2H?�Z��w3�=m[?R���H��^�7R�8���f��iBRo�W�7"��5d<B4D6���hl��Q��[�"5��#n�G}��4��q	�9��/��g� 
6�1����3��eG�OĦdk�B��5i�!�\I�A*x��� �bAUf�O��]��]b���%'ɔ�7\#߱Q%�E�_�۟,�/�	Q障���ϑ����D��.X��h1��:��3�'O�6r�U���V،-e6\�7f3P���__�ʢ$𝙿_녅S��v��B�P��`�p��i�k&X̕6����*}l��.�;��N>�@�	��X#�����+�-���?�l�@�ⴛ�S���|�>�W+uWei�ʺ�w��CH���A�����"�8��롲k�@'Q1�,����9B�M�h*Eb�m�b_j�z������r;UⅤ���+�̫N�zP�F- �L5d+��UNi�������u�g,l�t#y�}����X!���<���>�LwIa��|7�_Q�L:T��?�%w�
��3y�G]����S����zb�����+`�[�;���m�9��nS��2j�Ϭi���u���'Z-mg���^�������Ýq���U��_B\w4؛�?M��g���r��I_�lAzj�\+��ň����9s�:{)�g���[T1_B��kt��ނ@�e󺟪o ����������.�~�T2B$���]�P`��Rl�.�=΍�\���=�R�b�ⴓ�>��?�;���^!�nν)Z�Ǚ
�6~��3�~Y�t�C���0 `�!���C��V�1�N�QL=KJ`ߕ�ߩg���������T��������<����9��?�D�"���0T����嗲��]a�r�-�@�2n��:��"m��~�uf}�rbn�1Ĳ�������1~��n	YT	9A���x�3Z�	ث����O�V"`���`��C���$�������(�q$Р��@*���Rpk%�i�e�Iw~�ϳ�4(�/Mpޗ �8��8�-dU���ß�F��2U�t_ƋeS���t�HB��#:�Q�/��~��/�u �h�����I�nvT=���g��m1O���4Z[՚�A-�)�>���>i�ԥ6\"�Ni��s>u6��� ��u��-ՠ��1���o�Hl���>���=1�ΰY�V@���D/?���F�c��~H�+�6gy���u<-���&���Q1�a�Ѳ�%��A���˭��Z^�i@7Hujf�?6��[�u3�\�M!�I}@�6CV�n�,��	�K��\L�V�������b6�F�W�B5�<�0ƽ̶ƨ���vQ������A�v���d�*�G��ǚM�8��K�j�8Y��wIhf�H^pc�����w�{��?iG����٫%~jV��K�Ɖs�*�	�C�慊&�e٧�U>*pF("'�n���C/+�����_JN� �?���sFX�%�}7!TK�w���:�08�b��m�X�AԳW�	���A,�� ���w�Q�VG{���_>��*�R���M��q{�|Ҟoyž���r);8�� ��Q��z퉛3�4ͩ�t�b,qs���,�g0j���f`.MO��:!�G`e���4D����`�v�0v,+��i�����
D�Պ�ݚo�L1Y�d��Q_��(a+��̍8A�/e��=��/<*]?�O�y뚢H%wr�O�U�����{�E�c�jX����y���騇6"��1�� ����Up��+�aș��&��m�2�����D/1�0j8����i�q~(�RҒ؈N�ĤM�������a�NfLÞ-H�|��V$��j�<��b ��z N9�J����V�n�]��?���^��M���1,�7�u3#R��'��꣡�"l��.�SwoB�g�Cs�d:n�R���x6�Z�[]�!�P[��O�őb�v�ׁ�!�N�m����DH/�U?�f�2K�P��@�yeP���oK��[9�"���cy��V�
��xU��1ǯ���N\��"I�H��&9�EA*R`W�_ӛ�d�Ͷ�G3%�I�V�
B>b��SӸ.c��x$�Gi�$�#����ӭ���.^�7{���Z�9�W0���RL����zȰb�R�$#�:*+�N9[������,�t,-��py�Zy��}#��;�$d�~=i;��]�*�x��+���ī�*�g�o3c�����>�3��o�	` �N<��!!��	'a����܂�6�/����]���~L+4k!�*I�v��;��n������/�]_\�����H�Ɣr��^-?��^l�n�ܸ=8�r����@t!H!Ɗ��h@��c�qD�_"��s�����\���T�0c+����ǉڧ���i�Ș=�9c͹i�ǜ�����j�Y�(�ϛ��������h[�,��,���|��o5�ٙ_8? �Հ@��p��W�T�>��n|��ҭ��F��Y�Ґ[םma�| �� cX�at�nsXBH�M�<'H����iH���sL%iŉU��s�BoJ�E�|Hp����Or�d\��X,�C+𥳐~����B���vV�����ީ֡CP�W(�a��g �Fb-J�~mc�� �k��L�l�Fh�5T���k�S�6e�����<�r�։'	�m>��ډ�mvX���G�s�3<+��!�X({k��E��Ғ��%��b%I��������q��(������V"<��Wd�q>M���r���ձ��q�~Y����O��E���<�:~7����H.�m7�|�.�0�z�(�w�B?sW퍙%�a��
-�?u�����B��&p�7��I4t��kO$%�:i����kR�h�i���tP��1�)ȆO_!�!E��$yײ���k{\70m�-Z �	m�ԬR�A�ЍK�)ŉu1Fw�0�f�	y�.e4�7y�d�&|AU�p�����Me���Ȃ��i%~�ߞu���f��-��������Y���K����ۭ
�>�X-Ȭ��xq�f.<�Q�D�V?�'�l����ڐ��k֣e4At���Q~I�]��Ҏ�M;�Ӟ%�!�h_t/Q8De�v�v�/W�nۀ_ Ȇ� 0~�|�ʦ'��b�Q�G�tս�Ћ�y���t˖��.���|C0k�VK}�A�������a��2�=0�.���L[k� �R�
9R�,��׭ߨQ�G��ސ�e���f�I�1�K;����` Ҫ^����;�}� ��t�UJ����U��жZ,���<���OFhv�x�	nN0 S�řmT��~�	*T��gyT]���'E�w�\��d2w�h��`�9mJV9Xϸ5뫔����?�&'�z��
!ղ�=��TY�Q�l�c$Q.�^���=/E7
R`���B7n�c���h�X��yȈ����_��N�B�h���k�/)��}2K�k�+��s����H�լ�J�lu�(�!��ÔSYE�$�3g�[���]�#�^9�O���`k�p����u�3���_��&����պM���.���$sT�S �����׾ɀ�����F��@6�V�t����B��\��?����@`�� o �+Fy�]7�b��7�?��<b��_Wj#���Rޕ�y��c���R��:�08�[ ���H"������j����U�~�/���a�;��n�������������9 -wm>�h�>M"Ek�CAxd���#��@�밐���!(�X �S���Fu-�� �H�V-G�g��K����s�v?�]Z���Z�`!H��n⩟�l�slZ���$��*9��|�2�`z�o�0���!��(�|b�N��A U���2���`p��g�����F�֠7+oM�IR��N!R2b�qa f���~�N���Q��'���S�+p�>��R�
�b+��k!J�_��'�B��'K&�/Vzk��
(�j�p�(�N�	;����c�M���F��������h��yAe�]^H�.'>�`��XV�j���1�׵"�
hv(M��O%��,���;JH�3+<iҕB�ȭ�aӖ:�/��y}��-g������gZ��9\���C�D:R�*�v+��2js5]�s�c�uu�_Q��40�� +�7�r�i��ac�N��+6�:�h&�Y��Y�� �	�=ݽE��	�͓�ױp�ـ)C���Uy�*@�G��?�a	"ŋ�ݫ'١6�m����>���8RIy�h=�k�A�O��hAbj6&��;�)An�Ռ2u�������Ԉ�^�OSs�hFM�B~7N�4��p�Q�a޾��-�م�Nl�@V�A�8f�G��,�h��۽�2�yqST��^N�קB� ��J�|�T�Q�,�c�
�&�>+ߥ=1l�N�r�uEH���ڒ⍊Ҹ��]�W�B79�k.� \.É�.U��2
	_N�G�D-\�0��z'X����=55
UZb6-'�7�Y�q�����/��{/�������[�j@R�M��V��RP &��w��� 0KI�=�@>�1�,NJ��{�Ho�R�l�D�]90�
�q�qʇ�T]��L�ɺ�,��l�WcOlP��y��͝T��,�n0�u�l/NART�x�1`�[�ΙR�������Ái��WI�D���9����I�s���֐���=��S1��Ѝy1i
�P�量B��˾�ݚ�2�I��]ɨ߃���u�}���G����1�F�[���O�l�?�E��Z�)�Z�q��S��ڼ��c��@0�T�1�^}��'���Pb�Kfom��x�WK�ri��6i4�����ދ������dyE_�g�sRV�&�e��#?�#�Ok��$Z#-X�V�����<aZ�a@ZB�n�@��`�픑eP��q�ԯ�w� S�8�5�4���Q������Q�1����F��,�@��S�pT{�սd����y��?(�V�YmRsU���k�7?q5�R�-�V�.�0�>��A�"]��Ԋ��!��ъ@p�pC�o�&�2��t�*��W7w�E�v�'Y���4W[�kU�kL��a{� ��won�6d�{�7��0��x�:5���mC��>��`9��Ҕ>��mB|L�k�����UA�Wi�Q'
��K�W��a��Oߔ��³{���jg�`(9s=i�����F�h�X
�S�H}*������9�dI�m�<=�Ԕx\�:<(��z*5��F�\͍��lQ����*@s���y
���#[݀O=��h�Zӕ�E���ao�m2g��8SߢSJ?I���Up����������+�R���C�Ј�p7�Pѭ�UZ��J����&�3�d�Z�u.�*e<�
��X��Ŏs`��)���ar�i�z�N��Q� v�T�u3]M�Tx).�&��g�
U}Ylz��CrwW�AHQ	=�8�.�6��M�
9 ��ح��4�����;�$ʊ�z�<U�eS>(�/��"�G���˙}��a�+z������PL�?$=x�vG�c��r���d�����_^���������&��b�92�KL�4m��j�V �<������%�-�v���}��s��h���T��U�D3-�(NB;����}�Il�D�w�
4�l��� <\Dͫ,�W�!���+!�R`se?�����:o�,\�Ɛ�'�I�<�_jo:h9��˰8���E.��������"L�����p`����X�~I�äJ�'�H^;�+&G52�l�w�����
{�i�k#�w�+c<��O0M��_&{���FEU�:�H����M�""]އ�
#՞
�H�RF�a�td��T(N�idՅ�x �J]@��t~�unۘT��$a����n1[�'�`�p`n�[~�����؆fD��]�ٺNE���d�b�Y��ڊ�5�Ò~�� ����C��,� F%{q��!<|p�$����̮�pm�lsM�6�Ep����IlI��w�e��gq8�9�K4���`�&B}ȳ�em)]�1+X`*�e�#J ;�`�8X����N���<o�=�%W2b�*��_����Pm9}��4��"y�����Vt;�2
�9)��k�����2����<��3h쁼^30���R4 ?d���"X�_���|�����=ȩX��^�Y/w���}���.�@[�G�/Fݱr�z����ާS��K�X������UU�	�O���(�a�3�rarҡ�wM����-��ܷ��*��`2xQE%|L���V1�͊��Q�*�VD ��m�����N~����L�{Ϸ�Ǉ8��5���K��cڃ
_)��~�;M��_dΏ�s3�҂V�ν6�sϋ������4�
}��n:�5��'�j�zd9�Y�q�f8�C���SCw�[g"64�*\:̆�G�4��1�ϲxI����1H�k�\+��Ay؞���U�P�������nAwʏ�$�]����/�ϻQEJ�)�Ǿ�k>��cdp0�X$���"�{�]�51DE���N����Mr��=n] ����7�;`�G+.yYxN�D��`v��r��%�9��OVRN�"��`��Þ���')�'��O�q��E����<{e����ս�W��E̷�
��e�,����h��煂��M�N����E_�;�w���=5�m��k�Q��!c�z~I"�'B��܅Q�����wYc:M��1c�S^%M�������\/ݤ�N����c)5��HOQLI�i�-hj*i�NC�&����MB6�1�������Ϥ[.`���m̛z-��������!KK@�����U���q�6颮�;ڼ�z݄G]A�+a�팁���!(���Ÿ�="�\��*�����dp����=�'��.+��׷�=v<�y�	�4��l�^ۘ`��DԞ���sC�{�*;�Q���Zcsƺ���<9�4���>�I{q�k���ه�t����:�j�!��i�b^Q�9�\���S:�Dܺ|�
\�H�k%�����#�*ɫ
��!�we��v��{$<p����g���kn �1�k5#l숎���A
�8"�
9"nE!�����EX�]�.Q������P��#���7�(\�ךs.uh�xyp�v�
�l-8-7�E�P�gi���QG/P�#��ewR����J��la�.I�����.��~ph��DX�lQ���)�=�6���Xy����!3��=�(p�Y�K���=�%߆�(�!6�I��	%[�Ʌ�����t+�}adf�D����ðc�x�Ǯc�n?Gc�{n����@2�뙢M�_ը�l�{�q0ڼZi�G� rbx��B�V��ZW��nd� �:l��S{��\�'ҩh���ڿ{C��S�@�b�"W�!����42Ɂy��T'�č�e�@�s��Ƈ`���FDHl�p�c������/�^��TH������o�Ѳ� ����ﲖ1Em�ؾkgh�a�)2G����)��n*�H@�C"�j��{i%z�/�{ �f�=�ql��������k�.Y`׮D��J��H��/���y�\�h��O�y�(���� ����=�5r���Ƿ�	&�w��+�)�>����H"r���(�s���-��н��W����$[�r����~PTӥl��G�_Y�B�nft���ؔFOq�#�.�f.�s���R'<���yH-�g~Sr��p|�&󿍷W��Qx/�6��Ë���y�D�t6�jp����M&s����|��Ǯ��f_����~��)��7�/�V��@	�B}��wI���d��tz���4�^�(D�6��~��LՖ��gf9zm�'��E=��F��wovN��1�bK_�s��q��o�*�E��,��GZ�%*]Wu�Q9y����v��w4U&w��6:��q;���F�'ԩj�"؉u���MFE^� 4����C�����Z<#�ulQ�m��h��o_��7>���cƔ����k�*�;�Ȥ�.�iD$Zʴ�b�f���߸ێa9�F�b�#{�G�'��	�?R1����@�z�e��DD�n-P:�}m�[N�l1��XV���;��K��;�NrqږU�ԧ�ϣl#�
��C��y�:Wp�l�t����E2g�*'�+�{�s��f�(���jX��vR/�_��*��5VL��z�����B���������ّL_=Ij�d��{�ݷ4HQ2�g��w�i�,S<�p���K��5%�x�,�4��rdM�����@t���
LRI\��y���Rmݩ��< ��PS�����)?�p,Z{$�����/D�$�_�xA�V�����O�O���E�����&����Z�{/O=dw�N,4f� �A�u���w��(�P��UChg�M����Z"��m�Q�����-,��{/�{�����D{��������∖�¡bn��F���~�(�k�X^b���';?�=�[u�G�J����T��Z=��,�F�t���%�,DB3�ۗ�n�l�W:"�=��'r�3�oؑF�"M4rG�:��0,Tj�D?a�������Fo]���"��~R\`����+.�u�,g�.��w��^q?S� �R�)�ߣ�f�<�o�O����Y�Y��y�[A�q��G���jn�f\�k��!W0M�ǲk���R�hb��������b�,�,~����[�/T�����Z�UG�O�<���Cz���틒�R��G�����v�hĖ�37�]]��촒���W���nkusY�lU��qlE���.��h�ב�����O۞�Y���:5��KA�QK�&K�ϐϡcF��~����"�TQ0�h�dZN���qC{�cI�V�v&z���F������5�,L|�G�Υ�o� p]�Zvg�K��SC�C6+^����o93��p��ߔ�xF	�Co�.ZX֎Ϩ����j�u�;�(9X�fYNC���^S�� `3;y:�%�E^v[��".V11�ʪۗx�o�G�����������(H3�4��O^f)h�}���"s�]B���1ׂ�"~�
0i��˲��Nxd߼	tգdq.��&#�ߥm���h��Bד+�Z\�5&��+�]nD!Y�4ߔ�ܣ�6-����-,C�QǽB�}��j)��m!'ש:�ǋ�A��Ųa8Ϸ�{ݳ-�>��+���!��Z�g��۴_"�������N�xP� �n�ë<lk�VǓnćy+�R&�Y��/b7k8�5��@��HN+���T�H����4��K�����Z�'~�bﬥ@(f?ֶ�>�N�̠..��z}#@.�H��~l��%�
b�~�� �bЬ�d�굤ɷP�'0��I�c�Q��ߥW
� -�U<�l�c�x{��S�.�mwK48i�!���[1'���bK�d�⊏<˅}����5�"ǆ4HV%}�7˚��e\�:�Z�eg�*{>��eu#*h=����c~�W�A7n�ӎ�#̍)��1Ҽ�M�YR�I.�λC�Y�<��+} 9�h�'GjH_�q�4We���&�{�e�n�9��w[�p��l�s+�˿Jr��Bv4���bR��?�P1i���Ge87�`�Dgr�.�`!������0Y��F���&a�e0�B�}�po�?i9Tpʎ��=+����p���C��Y�!A`��T?1t<�4 �C<��3&��ż����ǛL��4���~�^�.���n~	��F�35�.4�>�г��B �]
�_�gQ�%��a�Ja�ͯ� QCk�`\�;~l]3������}��>Z3��F,�DF�&\�,���5/u���Uw��$�?j���g�.���F�3e� ���M ���+�Da/���Œnk�2��{m$H��ϊ����) �K$t^b%"�C}���Q�+7�I����h<��N��`�H�g��qP�(1_�������*}Xt�s&��ZK��7���v��� j+�Q�[�hϣ~k�0H��x�FލE�1������5��{����F*��H��] ����>S͒��i�D�k$��t��@�;����
�fNP?ȱQ�C�F�jaS��8�|E��Vm�X���n��B:m:F���N�W�N���EW>G�������� ����ɗi
�=������E�����fRo�	��oTO�`"��ȶ���&<\'Г�]���G�D�|�~��7�5�=П�NK`ϸj�n��(b`��?D_��j�>D��۲��XN'3e�_HF�lu������`
xL=������T�����:�g��jqڇ�+e��߾ZR�4~�E�9�C�}�)x(�?�_��3!��t���	K��w�����[��;��'��1,#�����>I4dd�G�-W�ʇ�o7R�7ň���R����i�ם�UN*�I<���9 �hy�ͅQqc񬤣��!��wi1C�0��B�B{4LH���$���╵ܿ�c�v�������_�~H}I�ݿk/��R>-sg"�a�F?S�&�I�{t_�Ԭ���_յM���s��6�����o�k�y�6���K	�;��7����Yre����@�i���A�Gg�0��f��cI5�}K�D��f�D����� H�2��dL	�����'��uN�hKh곷�\� ?n��ä!����C��gr�Q������2������t�N�^P���>������YAf��A%-r6����yt8�/3�I}��n<��+�5b������ e�����/cTyٚ*���6w/w�0�*��xg�A���nY��:��߯��s�B�6��&���*��}<����9��D��Pv���J�h�K[h�x6UKk⸛��/E�{���)�o��X`'Fނu�İ�{��4&~�f���M��Դ�-�г�����D��[�cg��N\=�?�t��?��;���Ы��k�wT����:0PQ�x0�B�
�s6�9�G^�P�H��[��e���N�F;��>��:oW:�����7àܝ/5B��+U�BY��>�[^�ډy���'���X=���@6��� H�)�X��5u�CO��7�3�V�����1b�l�z�Ӷ��ъ�P�zVKVn��|���y�[�>"��V*�A^ѱ=/�����b:��Ĺ9&Uy��º�ʺ�nz�j�2�>�3b%�շ�}y̴����j��"�2,�<�LMc��7ą�J�l�ƪY��W#~(X��j+�*7�)�k�	ɦ~�Yh�����,��a��ŜWq��x�9�}�W�0G��h��%��5�U��@5��u����y��t�"r7%��R���CH9��^�bѶhr���F�tN�����Ԑ��!�WZ�wLM/�F�zjK����z�)�d����ލsq�V���.� 1bp��� ��m�O��}�
��j���`����'U8��b���(�t�*���K�	i0������Y<M�gsr�H�i�w<id�ص���rY�_�0M��3M���ͼ�AON'�`=�b�d8A��'"}����$} C�ǻ;S9ng�?e�q>�n��7�U���8���9��ð��L`��g�X�c]>)
��z�ħ�]���y6��26��I��4��A׊�����o�O���dU��SB�ͷL�,��I�E�:�O؟=��n��+ 6O�>�h�,S��EC��a2��P�D��/!��fL����k�ϏZ�Lu������뙇.DF��D=����`����w3��S1P0i�q��2VX�uӁ�b��rW�ci�$��o[����X��ץ���x׏��J �yw��T^�j�Zc�V��O<�
?��*�yA��/��jK/�~�a���x vH�o��T���{���oiy��4C�O�S�O�ۡj��j�s�sɔ��π����Qs�t�C�e�{W�dX���F�=
G�3O���6��S"5����*����J���ٟ��Am^�{�Q;���[�Yg�@���D	�%ļČ*�����ؿw���,:}�8�9ƹ�ahQ�$o��=.��L���z�6��%,�Ͷ��7K��<���2(9>]�)p���ܧ�~�D��AO/�Ds./猋��P��S.��P����Cs
����Su�և���FrG��B�� ������c�%ɺ-��H�������S�<�X>�7����erI��?�a�N3$�]�%������bR�G���I~X��\&Qj8^J��wF���\C�� #k0��>��|���|�������k��e����^dKDI�N�c����f`q�5���[#C�ʮ*�5s��l��G�F5�/�<������p����k~5���
�K����>�5�WF��t�rm��R��g̃J��"r^`ig��U[ԓ�*�Co-ROg����Ч
cɹӬ�<�p�vw�1�ۈ���a�� cº��w����>�R��o����l`�-�P:	�L}"�-W1�O����n9���4��U�\@Ӌ�7�]�Bq8>��!�ɔ�@B��e�#��Ȑ�0��
�En�H�$/���=�Q���sS�a_�熋�;��\@(��ɴ�����t��iN�)�59{��v����E���,P����A$5$654�f#�Q��Yp ƺ�;��W�6cl��T�<���W����ص) ��t�J�2k8�1_��G%�ݬP<���-R�%�T.j�}��C�i�g��IiA�[��c#��w/���J�9�����^Jճ)��"�����˶%��QJ!B�j"n[������Ȭ8' >�񉐉����e�kW�W�1d@>p i.-Eg��s���_�s6eҚؾ$�a=h���.�R�i�t�m��A�x��7�Ӝ봝�1r��ٹ�zmJ.���)���#pw��长�� ���K7uMc�A}��o�ل��!�
p�<�)��m�"�2::5ܟ�y�iL@:�qh}_7�;�*��Y`Nպ���*F��@~����#\ِ�x���4�y��=� ��nw�8�t�����4���AL+��;�q�*���/lZy�2ꏱ�"�BO�2{1�t��f��	y���wÜ�LSr�+��q�b��J�F��5a�(v)Z��X5_D�Ώ�����n�q�Y�3SU��~�c��dT�wwFTSPJKrޓ+"_qrR��s|������ة}e����@?8���ߘ�o"T��\�!�����p����a򡤜���UB���,G����Mf�v(�$�K��oפ��Ň,	F^s>w��La=�露��
ע[��_�Z�������^W&7���+��mc�$7��7�I���[�7|1���ێ� �[�����$q7�D�58Y+��Xa}�5��A��K��(ٲ 3�m0a��>NF|�?����DD9�G�$� ��� ���������u��)��e$�l�����My�@ ���a�9� B<�~]�'�'T�	u
���|�w��d�s"���UՏ�vO�"t^��Y���6���3�o����������U�?}�B[9�G����*���(]������6ө��	Cf�\���|uXt����D�z��#,��cB/�D~�UcE���Suw�������
x��?N��U+,��qR�hK0}�?\�蝾�27�\u2mA��_�
�we�#��c�U�}�R��/��P���-�f�Ѹ��ð��[��R���%V�쥓�$i)���"�����鹰����6��%F�H��\��miX:��~ڦ��)2�Z��e�T����n1��D�<�UId��L�Ȁ������x;oZ@z0p�3�%�za3N͸��<u��3��|�E,A�iH�7⧆����9�����b
�\���'Vh�oC�TN�za�
bcPK�ofe`Q��.Ox�b�w(]�Y߅f�=���9=�۰{��
}�)��A�G�8���cf쪋�Z�Rs1pz$+��ۧ��d��m["`tԞ�t$LN���쨦�:N�L���&����7�˥��tz}VBH�^�'06���휚 �ޱ���]���o�"�E�$��f�ᴆ�W���8�H�s���|਑&U�[s�>���ɏ2����p6�a�NE`��>ɲ���T]�aw�4�I�0���p1���e��}o3�
��0�n2��$����&�aU�^n,��PB��rc`8R�p�TP��c�����?P^����ʂ����E20Y
$��<o[A��۠Lض?��XpZ�(�ԫyc[�e؍�4���G�B��}\O�\�ձÎҤ�`���d����C�%����d�Na��t�(����'C�a����^D���+T�Vĩ �`_5�[r櫗q�����}4[R��|h�N�JQ�զ0�wF�`��AV�sԋN�4�3��/��9O;�x�@9�_2��7Rn����iu��7=���g;�-��Ǣy���( s4���K�҄k��"�>g�������\Ii[�[{ox(0�����ZI���}e��f��S>EPC�����w8h�X�.P���e#&�a�($��.��N._�H]�v\ly��9����0���ba�]Jq6ߥ�u��uDNA�������и�5E���-;e>��7܍Y)��2}H�^t-U\H��]��.���(�ᶵkj"��\�U�]��k�����˹L�-�] ߫���EC�-K�������.8�oG�H�b)W�̼��Ϻ�4�'�� 
���t�CYL?[�� �+^ k�	��5�[5Z�TNX���k�#��n�}ͧ�����昊���A���tɢ9����;x�8ow1䯈�<���i�����*]�rO��T9��0�÷�D͈���S�,���rv�����/o�f0+�����C�����ú����0/�oXwd���.�h�W�Ը)5Jrz��A��#��mQ��:�[/oN0,&��PL�U@�3_�j���$�"qd=�A�9A�R;)��d�n�gk��nI޼HU���L�6��<�����TAVc㷱$���C1�hx7լS
�NE�x%��������Ư�ۉ�,�����{���O�co�U�B\�VNt������8��!&��4AT>���^!���L�4^m%B)��<@��,��]�4
ZEc�e4����(+��{W�@Z�e�-�W�.�T!b�&�\�Ꞡ�t�7�s���N\��Z�	-]2��p���4A���w*���:+�cn�h)��#������+�0�J(�7�S�p�� ����'���ό����T�U�.1�V>�{h���?q�Y�������w�V	��e�QՌ�����YbQ���|8��)ion޹4���,<����g{d5X�WLM&��ڷ@��V�a?S����%CZ��T����.����A
��uc$`19��V�S��#�,6�s�:HBTȬ�m�QR	�N��-��(���՗=\������cbJ���[���M��y+כ��wA�a�\|$0#�ua[���FԣZo�9�*�W�P���Ǣ���ʗ�5�Fn
�szcj�����־�f��]�9���Q���-m��Yʹ���Y��y�B$��	�u6 V:[%��II�?h0cW������8P"�ixWGr1���b3|��@�1a<�Ȃc���t�=�
�6�~�t[?DQ��Hr���2t蚊�g@�J��Z�[�����	�����q0�}�L'R�t.7f�$K��"2�Ը(."��Јwj/n��r�l����hI��PR��뤔o�6�d�T��R!h|k��6No�&.��D���4�K���h'��a�o.�nJ̐#>F�B�e�g-�TMAk��&Ʃ�#��D�7�����7d��^g���A��t+ДNz�EA�\VL���� -�;2�Nt:�=���!c��J]��h�!�6:8�`�����me
�W�u�j�g
��9�~�^{�oa���V��z�VJ��2��$� 3)w���N�\Q8� �7M�͂|9�{����UM���]<��3�of�!6��}K�6j˽�b�f�n�Va����rSE��wfi�`�����a����-�L���<��|ÌG񰹤fΘ�#�V\�wUy>g��u&C-�ʦFE�F�����$-R^O�B®Q��Wo�%%��ڿ;wgcgF��&���X&�Ԓj0��`.��_/%.Ga6�cA-���\j�*�g9@dv[���>�fe���VƲڮ�Qw*�;��_V,N%�D���p�%ZtV�宀~BA����Q���*���F��fcr��8����=�uզX��l�N`������/�l���]e�=]lq_
ڿ�R�������m�+qЧ^��S�?�=V
b!n�M��!��t��>N���#�E���qtT�m۲D�����N3u��r�\>�;�bO�1�����-��E�a� {�L|1;���We����Sx�ri��7�bA�"�^�.ᇫ.�n�Ξ���B��%d�N��
K��s�\�����D��`Zc���Jx��+u5(�V#z��c@�ro���u$P�������yW�\3��Poz"'XDf�
�f�:�:]��7X��d��
��~�E��/˚��5�~�?2�LR4�J���$1��� ������Na��VT�h4D��J؜&�3H���Pͮ��Z�Q"6��'ꍖ�t+S5
u�6���΍(�q0ʶ�R�j�H1�)7�y/���"q����I�ȗ��Z@��E�15顼��ѭ���E�1�0 ����N�8� ����?P��o�;t+�fV�e�qv�;Cޑ��۟	�������nz7\KK�;���Z�����/�2�!�:�Hfꔇs�@��6��wgC���l�b�����6�R���z���r��si�ߪQ�`ͮ�`�	�L��Z%P�z�j���Qoڌ$��s�l�z�.�6<�4�;1���f������Tɕf`WejlS D0�J�et�ڎ���n�i��#�0'+;ڎ{K�����7�T�wNl+��BY+_�j�
�h<r�p�X	����=\����.r��[O?���p���7�wYa�<����4l�g�%�o��-��p��z��Ms{~��7V�y��2ً|gY��o���+�ڪ��%�޷6�p�����C}e;���vk����.�Q]��u����%� Fl��d�uG�_I%%ȕʋR��{�K�{�η�H�QS���'�!�d/޷�	�Q��k�c�uϝ-iH�|�4A���ڷb���ӻ�h����n����<;���}L\�v\��i� �Q�����CJ@�d9Z
�n�h�7�IDU�Y(��-���k�r��{k�)��:�͒����d�ܷ�<�1��)|h"+�/Z�uFdU�;��轴�aU7P"0��%�%�aΑ�@��^��Q� {%G��J�9QH��lJG]���SN��2p���z�I�tcҴQ,6���>E�����_�;G��`�o��gx�E@F��_����<0��[(LU�!m�D���v����Y��{#�]�!�<���e�j�[F�F�h9W2����fơ��]B�����th��3�łA�>Gr�+L'\�I"/iDt�(w��ip&x�=�.�?��rMƂ�lFD�6A,��w�����K �>
��+�x��IX2uR4�3�T!���9���QI71�k&��Y��"���h�խ�����o��`H�!�G�-f}�qe̟�4b?N���4���7*�rH�ёH��*'A���¬_P�������A����� �f�)����ׯ��`jz�k�=q��V*ͺ���4R�y��=��GХQ�ġx�d�P����O�$�e֝��HDye���ߟv>�盩�I�Ţ́�a�=�����E��|�?3yBC$('��*x2��v�V���,���
��<`>=��d�r�8�sݳEza�J�Z�'·8�g�h��(Z��K�?� gV��x�f���^�@l���N�&�NLHO�O6d�c�s�VW��� ��i� �� w�R���-l*V�A�t��z����-��=�Q�܆�bv<�t^�߿�I�-z�~���9�C�Vo�����֊��Ix��Uc�K��NG�S*�(ݒk��%�T�m�}^؛g�R��FM�\�:����퉜�9��ܢH�5V�yF�04������{1-γ_ӃD�:i��Ei_�׷�SGCS���;�].u"`�c����o��V�[@6l���֢���r�uIMGz�?TR�����������������M�|��w:�)aJܓ��E�B�퉍��W��D��T<[��1MS�
t>���� c����7��18��ρ��q���x���n�}�����Wzf�Ǿ��W"o���t�>����].EH�b��8`��7�sZ��e�qE�Ж%��1�����Q*�Ǜ��Ԣ�'0��tZ[����5����6���!S�eGBH�,�[´��5%A��q��J�w���~�D^�ҿ|��4e#��Y|�:';׷fbS�C�5m��!T�����y�@��&h�d�e����'e2�L�F(R�)v�ѽ���5܇��:������R�P�?D�u��M��u�QF$GR�� 2�}�Y��y���[;�,Z���u[���/z��Rp*�GI��4W��bN1��	URZX`zt��TY3~O&B�J��u�7H�ыm6�w�b!�/�`>�>lYN"�i3|\���h9*�@!T��8��e�H�f�?�:@����g��V�x-ӫu�1��g��WE�'g-Ք.���4ʩcěr	����mP��E�#�0��9y�#�������=<���žu�K�^�
'�O�{ڂ���	.�vǢ����\�NR�'���/k��"����6/�Ķ�ӫ& ���2�����ޤ��%V�<L�O^��*`s=���ڜel�<�c�W���8�=�n�˳йˣD;$���11D����zp����^�j~Ɂy�����90�ʲ���j��Lh�N�obM�$��,�[~��g1��c�r�9
` 5��!�tb�elN�S�������>h��_#�c#����b�چ����e�Rݮ�)UȂ����0�6$��+0j�_a�B@~�TBg��-P��qww�X� ;�V��H���G��&�F���@��k�<�R��J����.�1Ә!�����k��FK�ؑ|���q�$s�0�/�f�0x�������4� ML��^K�4���~�M� }"����I�uHp�w0%�{7s2*~���D�8j���]��Ղ��sk��p:9j��}� u��~;�p�gƺ��� r˰*��;n�i�pB5^�}���d��+ ��&d퓨\f�'�ל����lgٍogj�g��4B���)����-��ґ��<iT�O�ڦcߩ����45+�+)7��I�<n<�wu� ��/v�L� iaɏf,�Y�zܙ��Qnܔ�e�lI�
6�LVjk�ʦ)8Z&����>��Njٹ4!���]�5N���U�7q
���a0�d��w+���N%.9�~�"@�L̇! "8�v�L *}a��2�(�JvO�8������ 0H�M�q�+u��O�b�Z�Y����-e���+�C"�:x�Ჭ�MüUQ�=��L�Q�Ƀ ��P6�h������;���賀8�MV��K�}�Q��D�!2�XtT���_R��]�����h9��`(���E�r[)K���%��:�]:�I7���W]B_K�v=F��ٝ0��Lܘ�Z���|����?��}�1Ř�������C����	?���m����J�LY���n��v&~��*6gA��]$��d��܀5����eO���u���m�Éy��`�J������ҊNW2+^,����I�ov]�rF���CÎ����%@����aEne�+X?*��\?��:SG��`���cq��R�4�<���n5,�=ch�n���YA�k��8�A��Hz�f(  �HrF\,�39Q����M��"��i#9ށ%I�+C�Ǥ׍a�x)!yCeLJ�~������o+��d!Np��넉���g��7����{�4ܕ�ϰ��vv����%ͤ�3}�~�ug-��!i$���O�6�j�kXIax`���<�����_��� ��Lq�n�8K\4rG����@k4)�Ӏ�z��6��"ll��<S��2&�z�hV��	�O�~:�Odx��n��ĺ��5�އ����& Q���Uq)��SJ]îL�V3�t|@cmSSZ����YJk���e+���Wb�0�x@��I��w��L�Z��
��'rShX�q� �{��T)7 ��"�M��=�܄�EԘ��.A
�&��&.�(��t�9���}�jy��l2�de3���v�!�=78<P.�CX$�ӇI� Rg����F�*'w[Ux�	� ��ݏH駐쨻8�����.�׭U�B��ʣ�_'��A��n�O)��Һ��d�T�=�m �|���~�uI0'g�y�C��H�;�K���L�\�N�F������Ngp�9����s2�{G�q0u������_THeq�����/�h��ZtZ��Zl��6�P��j��!.dA��W���?��"p�+�����W@R���b�����1Ά�>�woN�لO%��΅s{��F���o�?��i=��~�G!%�$��s����(�j�W�7�q��k��0�*�2F��˱�g݌���q�$��Z���F�ؼ��O�jX�`G���b@$��fd�/�_��l��,�0��-��Gj�Ft�w�XA%t����襗�r]dm>!�W��3�kk]���E#)2����d����a˫G鞵�Jb�W�C���EH�j��R�<`]����\NM+���`��f K^u�� ��`�>A���d)?w�i��9�� ,�	�댂#�5�b������jع���[�R)TF���@	�_���O�9�	T���p%�`�m�a��ن(����On�(�t0܌��_�&UQ�������;�j����H����g蜵N;@M珫�6���9�.tzF
X��.�E�=��}��Y����R�z�`�=Q�:	Jgi�H	R�EǾ�@K��h������Mb+*�������m����jܟU\^�힢��[Q*���h+�� 0mm��oM�.��������D!no�jL� ﵉yaE����h'F&]O7})����'0��u5q%�|�η�0s��I�����c����Y0/���n㦤�|͚	 ��=\�5H��|�-%�VE��9���IP���x
�28ڒ�=�o3e�0)72C���W~BD�>S `�,�������yhs؝hǊγ\;�$O�J_�H�=�Nv��%>��L��\���l_�}���
f>)�f��^Nq�]�;"S:%�?�uf�2t�M���DOt�p��N���=�6���N��"�CR>j��
W�]�$P�s��EPj]u�1��D>��)i�_�qF�` Os_�}]X�j�H�G�M �xx��'5�
����,%a
6�w��N{��CYd���?�0�Xt�SQ񠉼��zS<�c4_�>������M��Dq�n�z˰��B��K>����V%doWT�%���>#���^�hv�J��=iI�Q�V�P#6y�*"�.T	c�(�q��%����Iq��|�BF��j&���x�Θ.��y0��¿s��#��śa��$M�0 x&��� X��H"���J;I!�����TTCr�Vٶ&C��a���$RJԤ_����pӧ�`�2X˒��iJ���]M�3��5n��)G��8�͎�� [��4�����:��eM@'���*Y�o�(QO%�Ğ	�Ji)�'�n�{����fl�ܭ���\ �SSv��u�Byr�ޥ?����� �^M�%noCٮM=��{>W+x���M�Ak���=[�K�m��Pd;�f�Ҵ���%A���?b</.:��x��D�@���峻�m��!@t��0HR-FaF���3�;0�|�)�2+��lk�9/ne[��T�b���ѮR�.�|A��˵��C���퍂
��bлb�+������\|��$v(��	������%"�e�M�`�r��Ǻ��.I�V6_�Z�ظo����6��A��l}�2��V������(L�D�6�dZʼ���Ȉmg�)?TS*�_	c�g
_�ӱ���)��H}�����@���ћ�����9J����������˳42x*�#z�+R�a5Gx1�9�l�ʧqO�)�<�*���Y�Ih ������@t�nGw�*�Y"2��^�R���[л*e�r�15��ب�Jd�/ )�oU�$� �`u�$j�/��4z��:�ᄼ\�7B|�6�&}ł>lEM�s4@�eQm4���#3��xۈ�y���Wro+g\Ÿ3>}G|@g
T�����Y�1s�+Tv����@wݼ~OWRa�@jV�;U���Ķ��O��e��@��h�
�^W#2�r�� =��hF��'#u��cz:6��8T���GU5p|����	m��}�ݬW��B{Z�M#`�!Db��� [�釟�u^]�cb�Z�z#��F�k�!��Sw]�^�f�{.��DI��u��ʆ��IV�vZ�o��+~AF�\���F�z3+�0��Ra��/]*��S�Z�v�Z_���X��5А��oC��t���/��O�	6��Y�t�����@�t�$7g<�J1����ș��T����afRX^���Ǹ^�������?�y��K�*���h��"�5�ƿ#[[�M������f���UF��!H�f�5C"YlF��B/��]#4�ƒz´�[���o�5��NT.�o�G0��'�1�64��;%։�ĺ��KO9��ųR��QsE����C%w�+ì
k<�{��
*��t���?��������!�]�pӐ�5�f�zgc+EfV�S���~��,��v1\ ��'��.�~r-���L��WN$Ɛ�(�aN��X��%og7�)�o�v�J�A=r+�)\5Q����>N��X�8T&�21*4Wj�
Hx[@>�5��H��RI#�#�)uO=����C�$�X��{���~��h�oee_�E�88K8F��c|���Kf��P{/W˂P<�|k������\{�P#�v�m˽G��X7g�%ʂ;5�$�"���؝��t
����m[���H����Ǿ��L�]��b$���Y �	9ϨT����A۴T}+����ևɝ	
'�U�m��S@���~|t%���g�꒹��aS_�e'W9!g������q������P�5tF���?͔�qʵ���un�)E]�h�y�cc��G��ɔ|��OY�Ъ����ʹ��>�O�J��"���1V��X�<��>@N��4�FTV(�ϼ\�<�0nZ'T�MC��gI�#!���Կ�#���.�ܱ�Z��1�w�=[�3S�-��"
fI)L���o�S�o��U��>2��zE5����}]�'��ϛ
�_���C&���r�#��S۾�(���^`��n�*{`V�8e��ye�bT����_ӴOR�.!�7��a�-��"g�'��{�q�&���^��-fpަ/�z�G��	��["HԹ����V:XC@&�:L�K�5� �GI�,2o�&�����y�΃�U}�n���Pg�^���_��l�f Xh�i�钂�r)���rI��	yRGa�U��"�SQ�֤����3H�}\����@��$o��RB�5t�"�&����͘���=��=��:�Q�ϲÚ�P���<�^^�|�E��T{T�}nKH�;KN��:�ݾ��e�s���h�Q_}c�7���� /-�	����~Q·��aP�Q^"S�~CJS������s/����v��~�� �(����w�s��_����|V�foU�l?�c�h�'n-�sd�h!i�2�!�4��U�_s1z�����V	�O���Vo��,ǅ��mw!��k�m�p����/ώ^���Ԧ���d����獓l�3��{��f��i,��hOW[������H��/Y�S]��DtS��'X�fa�U�>�/��Q�g�a��@�mV]P���-�V�~�k�t��w���
5�r7�3������F��=�lԋ9�۰0=�]y�=�#�\P4轥�.���}c��y�q�C�m�|2�+QyRS"φ�n^���5;��`Y���F��h�����lq�3�y����f=��!8�m�D��=���Q�lC@	�M�v%E�ˮ��J��C�M�lƷ�4�]T�Zr�  qH���f�],~UgLa�QP/5ǈ��v�����D�2�(��0[�QN(��L<'~S����Ey�>CnE�@��E�)�P)���c��2�[ A��?-�E�N�s�����m���n)�@A�z��	���֢A� R)�zP7tv-T����r�5*7QJd��5��A~<��œs��봪�HX+��e�zY��<�ϒ�q�>���e��-��D}.KJ���Q�.g%p���И���Z�����J�厒S���>������7��'�_kӈ
���h�"�9�­��ė2H�=0�3̉jP���0NW�8.������yM���\F|HwC��}�����5k���L� .�&�~3"�҂J@�TK��f��B�^+%}u�vji������ �OǊ����!u˹Mt�/���RT���s����k��fwY�kCqח&�G���!= '^��ؐ���=K�g�*������wP͈!�O�5��|� ��wC�*��aHSڶ��[m�A�'�O�/����;�Z_�P�*�3˗�FЅ�P�-	�#N�#�I�[�J?晭`Kw�B��#�+dԱ� �ǃ�VP����G!Xݭ�r�J�r}{1�2��Z*�1>Eִs��\����]��#�EbH=0;�b-���l��-��>���N���9�
�z�=ԛ@�q�琠�"�?��/�=��j_�����4m��>)G"���ћ�P(�Np_���^<�p�؞�8�g*Jp	
�>��ZK��B�1K��!�)�����F����W���wS�[��{��s��K� �߽I�4i�� Q����h�T��7�q:l^�"B���o)~�U�m������{�5/M,z$$��Y�F5�8�/��)��f�{�>?.���|�b �ҰG���cB��� �)�v�ܻ�ب�1�S�����B�K�şt#oeJ����"5��4*��� �zN�*��"����	�V�����Ms��{`�������κq��� M����`q�$�~]v����M�&���00����?����}�:���ي��aLG;��n`��3bD�{i��ҕé#�o��)��l�yZC�.q-K@�~pv�pڎ
�~���d��aZ�g�����b�
�k�'�D������$뼢���CsX�~�D������%[���j�4�n
]���R�X6�f�`Vt��&�����w�$x$j"�.�Т�3CI����_8�5��ː�5��Q�)��H��wiP�{ �B}�pDE������,��&Y*��_��rVRO�%D�\���bg��v�E��v�Mw�t
7��4M�/D�l�&�=�[A���
��J�/��׷Ňet�C�-iuYf�h�-~��Sxfwi�]��@U�/4�B~M��/$���-@��0��%l���l.�ṵ�;V�5V@�́6_h!m�Ȕ͛?o���l�~�p��%G���<do�� ���vH�i=�ߺ������[��Ď�!�f)_LP���/���C����^��]�G������Ӣ��9|��u{'B��M�һ)����H��a�!�͂�oCN�N��|��W䮟͡�?$�N�
��:�ŵ.���3���)��:���.	.�V��5_�I�Y�:����#.3�"��Y�N�c�_w���*V��`(C�hw��4�I���˚PdŽL���%�aW�n��
~�e�W�ϛ\�����4"��l���ن���eO-�ZH����聵W|��>0Z�H��Q&W�ۗ���߼�a����̭è��Y�;�(�8��_
ۮ�(f�ل�S�c��'90�D���G�N�j==Au�b���D��U�LS��x���X�R����'���K���[#�B�����i���������]n��)Iw,���t7�P��X����q��%���vI(0PSB��&z�
�E�~��y��c��1
HS�k��=v�|A�nk3��,��D
d�����ɵN�d�����&A�t��K$�,O\���ť��N���R����ǒ�;
��0�?�Q]�3%���W�9�����gN�u����#�lW@�����3��nUa&m
������(��'(�x~R���٪�1��t�~�}���&�tcw��&�p$��K�����O<"�mK�PRH'��F��MV�m�%�R����n����q�+"����SȦ���O����zy�t (�Y���G��'�L��6Q#»�����2{~�Iu�3Ց�=[N�B$����D��-��#�]UpS ���1P;"ݹ=6��?��r�yv�����2��ݰhGt�a��i`���;4H#��e���WF���wd���8�1�?'���z��_���Sݾ�e�Ltj0p����<� }7uK�D �D��0��_�ݣ��Jnn���ʇXWQ23�0�7��^/���"I)a|X�5n��T�j����?��F��C.1��U��F�'����g�AB�;8�i���I��Χ���h��d�y�0
V�l�����O��*��/,��=z@'�!�ѳ;n�(��)�I �+F�/&8��3���ЇG�PC�drXslLF��_j��f*ɪ���v���iCV��݈b�$S�v)�$��&ۢG��$������-��ϳdX�(�Kueb���	R�+^	 �0��ђ�Xj�DͶ���a�V�	(�'��3�ڜ�&��P��B�Gmx	��ͫ���_� ��f9���CCB�^�o�m�E?�"������K��|�V��a�z�e�ؽJ3Y�Q��5s�������N?p���q�ex(�n+tݯP�$��:�O��}(�����ۦ���	o�=�{��K-g��(r�!N��5W8�CbV�xf�P�s�<�e��#�X�0��\�����L��@�y1\����.�ż��۸('��[����J�h*���lbnb��e
�&�a�?+R3P�r��:��&�m�"�:�E������O��m�KX�nz�W���1%���	w"�s.[����pɇ6�Ķ���� ZS��?�}T+E�KH�`r⍷�����u��u���K���)��l�w��@�c	[sՎ���n��[�i+' �F�㺖Pd�QՋO��.�cM�����Ǭ˻8��H��%�� �Qm8"�� �i{T��rI�w(���?@���`
3��U�����z6�ș����{��߀q��M�!7���� �e"D���G�R���̲�-��?v�d��-�=�9�����Z��P�M����p*�T��,�B�5M6�p�|Lc�Tm�/�{%Á;��*k�W��������� ��7���(t�B���\I�eU�0eWT�kn�G˯��4^:���vx��os�r�P���:�IS�}���$�i_��wTI�Ӑ�n}�њD���t��n�N�Bm��ސp1;�m���-����EH,�]��{6|ٍ(��lj�^�K"[��G"F�2�=u�g�8m��51��-Q��R�����!On>@�V}�$��q1=�fQǡbH�S�w�3�F9v��/�H�����c�:,���dA���╸y��� 21��`���pB�u�(u+̒��w#��,F\.%݌;6Y��\��@@�N"��6 #~��Ke�.�b.����AKC/"l]��w�؃�!����䬅�6�^����yܨ�Ƶ�Il|!�d�Pݒ�����"IV�΋��!;ڦ�'/&��|�x���{"���#;N�t�vIa��ތɦ��FS�cE�3�Iѫā' ,��� a6�>u�> �_�'����l�VY�Zۯ�d�%�Z�XVD��/�����b�[�17�]�_��x7��Q'��r��y�9C��Q[*g|ǁb�"�F����ۮz�M��kT�������>�br���<�}���UE$K�]��^����a���("�h�'�a�y!�v9�L�P��9.N�&����_4h�#���`.�(�߶f�	3a�d����l� �f����ƈ���$*X��Zī�)e�C�D�+z�{�s�o�!�i�P���&�乭Vp�M�f[����Z|��a�d@"@5���,D��mp����p�w�*&ޭqx�\I���_�*�ŉ���"���,F�7Ht���w3��`?�l�H1���%��10��E�;�j9���0��FF��A2y�U=�w4�}e{^�W�v��G��6Z��龧�����Z�՛��ޠ.�쮑�FARݟ�U�$Rɪě�a��d��T\+�3�fr��$��Gǻtc���r��غ�B�z%��r|6�ݾK�c�#VϩLc)��	Ք����X1r��w�T̰��{%r�J	v3��k� [���y�Z�Xdg���}5�Z��=Ӥ��1�U���{%���؄g�G�J�6��\��{qB�󓹡,����r��c�cME;8�E��k,�?4#��͋Fa(1w��>�GzYv��HI���9�y�W�ͺ,z��������B���WU&&ѣ�o��BO�>p���A���Wi�]�o̒�8��j��׬���k�@���r�\K��-���}��^���!h\rzD�~r�T��ӱ�.O[=+�1��lʤ$TjP���!6��qՎ+aU�|�T��C��}���w�����Z����u���ϻ��PPQ�<����2���Q��)Tj���N�t�5�pHb��X�{ԟ˃xع��M�1jm�YI P��L��]�[�s�R�[���N�`��o�E���po�����E�)�ؘQ o��X���%Xz���V�)e�P������d<��Y+�/�}�k���|��CW��.*�#�^��p�_|�p�����1-�bDhe@�֛'EhgZ,)��֢8�;��m����1��ʬ��
��j�`Ɯc��!���o��GgNը��wΣ�)�`���������VH���0�S�w@��t=FhCi�Y[�Zn/X&�l�a����{���$�a�I�bb����	����d,t�p�+�&<��O�!>$v��i����8�ǎ����;~M�g�B=�H������h�a��B�/�:��l��Ƒ]
���#fh�n�',=���An5��'�@�오*�%�|596�EL$�45phߘ�CV�&��Ě�q�����9��ÈK�`��"�F��8s�����h>�����ۿo���~�Z�J�6+��7hj��0ZT,J��-
t-�_����qg>u45�1w�%@�j,�����H"�p?	��3�|�),�G�S������|�t��uEs^�.��6��\�Ɵ)��mut@�������}0�l��˕�N5D)$�SB|Y$��P�]-u�R���t��#�m�gf�5P�y���	c��ubw-��b;�>E��.�4��T��v��9#hh-��8�'��]T�O��])��@٫������'���9u
�?�>�������:�߬�?-���y/�Ň�t'�~r�ۓ�k�}�j�S�J�O� ����O��{�h�]�0A${�0YΖٛw��Z�s��K�.u�D2�j�x���5&Ⱒ�����4��y; ��Q�5)sO·͌P�^`h�Hc�z�+/���~��dԋ��I�a����͡j���6�*R���r$�6ǘ��U�p��*G
j�hs>�S�gc�6:��Su���'�C!r|�|�h&����V�l�L���z`�Fm���?��� ��q<ܰ?�ɦa�=�nT��k�ҟj��{�zOX>��Eq))�O���T�����
Z7�eP�a�tV���VE|��r���`Q� ��8@�|������7bd�����hZL&������f��U�t:>��ʨ��./
����0���ǲ��D���_;���
���.����ih�LIz��}N��Q���C���t��v��q�oC��p�*�N��D��u�M�:�ˊ�9/c����2�����"�K
9O�'���wP	����8dG��j*���Rj��������Ϻ�i������ ���X`$Wޙ��(�ȕ S6��yQ۹��8�L+�6
�E����6��Nl�x9��O+��x�����rG�%u0�*��&�Rt��c�����I�y�v��R�>���x�z�3r�M�u`�[<��ix��w���mp�X��#�l}ˉ��R���ӓ��5��� Բ>z�B٩(4�4BXT5'�Zi\�`���,/�*�N����wx4̵�"��?G��qT���&����N���.�%���&ծÂ���n��?]�Ƙ�=:n�Okp�G��K�@�A���K�
3�Q�t�x��,� Q���T���,;���y�� Q<j0����1�F�����0xw�Ge
֢�d�����w���g�kW1�y�;Q���(�Of�#���>kn���[��{͚�Y�z1��ۆ�P�]�:��d��
�ڥ\=B�aM&�ɂ�V$A��ɑ�|���/�h��;�a�^FMx��ț8?%�����O�1wM��rCG��Iu�F�b�����Y@��fv=��n[�#J+y�D!�GHqۖ�ȸ�`JS�:�H6�M�o��@'������x���\8^Cy�86�?cW<q��b7x1������ �h�]a���2JN+����c�Z�$�X�L��%�?<�I�SKć�x��&�X��^���D�]������E�U0[��b��{�EŅ��ͫ�)>,<����TE�|���n0�)�>��:ʧC�)�6(�El��!�{s�����w|CV!D����>Κଛ���4O��-�$�Ӽ/f=	�k(?�W�����o�����_ܓ�79�<%�E-p��.�c�C�=2`�������=w��>fS�s��'Rx�lf����@�6%�rK��|�9�牉-5XAW������w��Y������]NT\d��@���cO�6��iZ�ЃV�9d{j��{+������{ŢNް'�)�=$��#�}���"����Q������yL ����{�3H�e�o2�Ah��G���{�������� 꺵=�N���������c�t��7t�C*0=����3\w���d��C%|R#��:զŁ���!k2��	��=� 5��Ã}�p��+I#<L�����+���w�+����,S�0���D�h������*Z����<�B��_ݚ�\+�}�Y��NH�#��.�3k=�#�����jL��^�\j0��#eC+�E�Hj�M����Ц�1��A���	�no�MҠTͶ���sD�9�q3g��]BZ�S�EX×`��b�$J��˘M��*يc�'~dhA�ea�_�b⠝�^ǻ���@�I��������뀈u6m[be�N�|�ڿ��s��]�z�w�Z�u�������W�կ�De^�*©��^��yO\�М_S�+ǘ�5�=��k@ZZ��B��g4��΍6A��$8Z��c<�w�0v/�r`3/^|X�"�;*�zu��0�˓K�^aԙI}�EQ�[��GAhD�� �;���ĕը�P�����Y���=�_;=�	��q�|F�ހĠ�x�D�g�O�d��^ b��8J���&��N)#P��}Vڠ^mˮd��N�!������L]�{����Ɔt{r��PA�E��8��o�bAo�Poat5,&
G[�܋�����엶�v�jYe�T(NVF3�1o�G54�m�#@�>��66��LՔ&n�<�9���ToG*��P��l��C0��â\إ�'�t�荕-��s3��J�U����]좤f�󑭍K����jĻ��)�x����B�+�j���'��V�
 ����{��6:��+-�}:�k�ڇY������z9�D�aȠ�e��(u �6x�qUd������%�����"\�8�	��W��T{�Ա5B��P:�i�n���S��Vq�Q���m�ga�2Ć@V�ڝ���\�ι��-ۣ� g:��8�ٳ�Yh0\��0H�u���Z�X�MLc�V�<OP��z��S�7�9��8�b������Uv���<�~�O��Z�����ZV)��FGހukD)�A�%�ܩx7w�N8���D�����:��}
�j5�=��[R��sՁ10YeWQ�����dD�����t40�6�K(���O݋��A�������G�z�DP�e£�X�J5;H�������_�]��s�"�߳;�.ͥ�f��HO�j#�Q��I'U�zn�b�������֖�A���g��\L�d�&��?��؉7*>s��6o� )�)���lN5��������X�?���X�h++��������
�b�!���p|ם�Ss��e�����0�U�zbN�D9x�f�K& 0�8��s��Yx!Q�-[j5����6�v��!���!�E�l�s��U"�v�q[?ץ��b������T�t$L}ٌ��}9��/v�'�:���Jo�?*�e�~��c���1(w'�<b���W�u'�ǅ%�������߽�i:Q��C,K���Z����jY`�?q�ā샀���l�a?�厂�d�5ps�C�<*U�Z����2���y�����r0c��}~��<�mT�LD�}�7�g,Tt+�2j$]|� �n����w��w�^#g$i-��}x�(�Lp��B>�j���Tw�j~;ݕ챷^|<h�sY�(�-J3�����g�S>�D�-���j�����Գ���i#\�OZ��?�6�Ih(rr�J������K�]u�PV�P��U�q1i8@8�Fs�۲�E��JpO*��y5��ԏ��7bmVm�����<?���o�) 3��
�B�th����d���d)�
�eK
o@?�B�;G�h^�o<25˸��w�=K�A/;]Yrs9.����&���P$�����a�Mg��ig؛\���!��6rL�>�m���.>�*.�� @�B�N�R�0&�3gn'��WO��xP���o�js����TG1��a�t,�O�B��˽ �|-Q)�-�'���d6A �	k��Z���M=:���®9 u�/�_Gtn��:IWeP��i��̔Ԑ@�%�	Y5�Q��=8��#d%n�f(+���Ӷ4�	:y��{N7`�V�ދ�^�+l���%���ޭ�Һ!z�"�Cv�(w��62]~�_�ܯ��J��Ѭ儓����B��xa�`2��ٙQ��M�;��=ވg���F�[Y�\]�s;��8p-�5bA��\(rT����S3����ӵ�b#��_�?�P�����s�)�}x�dk8���;��ӂ��g���	~xn-$SK�:g�T�À���ֳL��پ��1!{s3w�֌�BX��l�f@�Y�1OWv�	�/��`]K4:��[�:�LV�fȑQ����2�V����O{e۟	��^����&��FQ�e�S6ޞ��Z�;T�9l��1��z���$���Py��J��疳βw�h�Z~g���9������g��H��l����@eI:��;�4��O���P���Q0*�.?�DI��4�)"61p<o'��E:�Gݾ���Hd	;�#R*��ʹ�J$�z
m��5�~Y���w���v)��Q�����SJ�F�n�^)OH;�C��DR�6-�I�i1�/@QM!����r�q}(�X��p@�L����w\�\H�0��ű���(��X�Y)��h�_r�r5䫈�aHRy��M���jF��a�����H�����:n�l�����@`��Q� %6�h�}�RHlכо�M��Z��|W�
؅C��-��X\��zO���"c�_pL�dUR�R�w���ڗS�P_� B�	v���$�=���uY�/7)V��	�;��Jh�3�^��%S���a������<�e�7�Wi	2`�|!+��>�����i��bp�$Y�?PC㪦!���9CPw< ���z�O�P���{��ĵU��妔?��v��?
a�_���D$�=H��cH�퇀��l%�(�t�j�|+ 2�KgV.:��2/H���h�o�V�| �Ull"�b���.Bű�mK(y0A���3#���o��bw#��7a�6fn�:�n�ȅ�,��p���Su,�����_F�:��A*C��!�tqbBE������$0.:7�n�Ò����h��&���Q���8׬�WU/��ʺ�ڸ��:v�V���U��wXU��M��Xt��$m`��N��7d`�^#��uȶ�ߓ���@�b"�Fv�K��� ��a0��@�>�~�����O]�ٮ\���%~�bˆ��\�i$Bt�Y�����/u�L�bRC�@)�ݛ��Ī-�=c�#� �lM�Xb2�dQ�6FxR�#�D�G��t+�Ve|�#Cku\E��+�$7.6�/M��R�^�dn{��LN��N/T(H��b���7��bF��Y��N���h�����pg���Ufe[f��pؤ�^��1b�������׀�2� ��FAd>D��� q�-
B�N&�[��z�\���skT!�g��~(�+�Q��Sz�nSa2X�÷���f�n�AŐՊ�e�5U����N����!w����e)��G�!��bU�&��X�V�]J��3D���JS�v9��"��?FG���M��g�Tb�A��XT�O�C�K�S�̃��{��h��v�6�cbd��#�xDW�8�ʯψC�1K��&R�/�Y�j-�-��3"��f&�`���T�C[@؏3� �!���~�q�s������Y9^b]`���BHA��D���\/�m&�?ުԋ+���v@� ~��2��Of�֚d�V��~�A�@��ʐ�͏��8�ɏ�x\HK:)�n,��N��_)#���6�	�[��n˚�5ĊB֬���s��jTq�U}3
r࿟�����U�c�%㽺D࿶;��Z�l��uV�4=7yN70\o|e��5�w�\rؖ�-�B�y�O��,n����D��
�y9�(޼ǫ�Y�M	�h�2+�iJ��NB隧?��txD9���o�Cj�l�.NJ6dN�F�(7uTf}��op=G?���F�0���2v<����M��r�w{nz][ �^�x��i鱇� N�A������r m�U�)Q�d��fG<��Woy���!%ܩj�h�>(al6^�u�7QN![pſƉ�(�2s�1���jwY#�ҷ�j1�+4��r)���i��*s�#�d;Ю�c���ڂ�x#h�`�� #^����!�.�P2���И=Y����nߨ�e�W���#;�bB���ȗ��;Z?C_G�C�D�e�A�g�%��,za�aŖ�����#H@yN���HrC����������.��!�x��} >0�cIF-��ةK��w"���j���zA}i�K�WKOи� �@��BTW�Z�D:l�oJQ\/Oi����բ��V�PT�2�7���G��@�5h�m�κ�Oc����(�ɭ�:���-��&� �t�o�n	K�"�w܃N�@,kwf���5��|����ԟ/�}�!�I�a�tn�,�f$=��y����)�/�>�. �rĐ
���N�<��a� i�s��w.�g��ؾ*[i�?����b3m�X�h.ҁ��Hе�V�W��-
�j���!��H.�p��E� ��1YC�����aTa�m���(2o���l��Ԛ�~R'i}Z�D����8��ݿk�Sb�hG*�,�G7�Vu(M�I��m���U����b����@��#uPue�:8�f�Q̖M	,�����+X�W���!�Vf��:ze�/�Y�~=�^U)��u���9�P0,ĳ5N���D8�+����l���r����r-��
�OA�:��wk���h��*�Ϟ.5�X	�~'��|=]��0��d�Le+lF_J�y�'���o��[��e/[p���Qܟ��T�%"�A��B1s
Ƽ�Y��j��ʆ;�8}�}H\��� ��*��7��i�]��5�w_m���K�#&}�?��]��Ό^���ߐ`�eރfK�+�sݡR\�����6X�!m8��1�e�Rg�L������kf�d=I�q��T(m�/��G���O2��^�݆9X�M�O�����>K��H�"�U5�`��4� �&j�}�HuGO�H9�9g�s�|d��)eid��R�v�k�]�j�$O|�I']C��� n��f���72�����Wk9+�|�F��c� tԽ�}���r�/1��'wkmp_�_�GT�捋�V��R���>�E��X���*<tPl��T��c�w��9b&�&�8E�{	�����l���>�_q��\����L��m�8k��F�腵0��j���/)��w\8��g�@���|�?3�Eu7�Օ���w�ye�^�z�kty��&O��i�ef�geZ�з��`��IkQ�{��;6�91�^����.��c�x�_���D_ QL��\���Qd��n�{Ѕ����Cօ1��*���Y�@;:tL��|����p���8ZB[����W[$�X(��X���������>�e�ʱزo�Zy�����K��@��-*�)�a>-�4o�!L1o����a�R ͮ��Ҡ�k��1��.�ݏ���]�rpb��F�4�W*��1�w�',\�̋�җ��t�v[(��~b��@p��j!�w�v���K	b�ܲ�DZ��|޼t�6�Z,��l#�B�V6���9�����0u:S�	�:G�e�ޟ�6b,�yS�8� ��2�u�w ��h>h���j�ȷ4`�,S���_�)w����.J���4M�*2��&^��
ɕ��	��τŕv�!V2Ne����s8"�ԩu1��PVlԳ-�*_`G�`��+������h�d�8Q�m�	uFs����Z-54�J�h�`��34��8{�c�~/c�����rA��Б�[�w/Lbq�x�#4+� eh���h ���0��`!Z11#h:��J�$h�z��pC�L�n��p�.sƻ���|��?ɺrY�/��G2�Â|�^N��)���9Y��g��pQ�
�K�Q�"�h�#�{��/o���7���@6OR347^:"V��;5ݪ=dX�ǁK������;��,�5�_��W\��<E�tM6�W�rL�N}E���]�c��,<�����mt�k�,�Of�Z�~�<Q�S��;4!>���	"O�5��g4����r������Vv2l�I<I��m� ��9��TP�q�W4��`UwĢ�R0����S��������m�X���]�I\��ɒ}�o�_2d�u�,�7%�u�Q�9Q\���־	��L�I��b0�>������ZK'��E1�������_`�����G	@&m�ɂuraO�����6�{۔��h[��'*K��"���Ro]�뭺�[qX�rޫ�$A�i�.D���y{!9��հE� $�vr�����@F��+��+�h]��i :�E���#-�7�G��ϣ.�bd麇�����)�@��*��nf:�d��Y6l� ]��5?zXZ��)��B�`���o��>T)߁��PU:�
j�>�`�M���!V�+�靇�u���Y%Ȟ���ǜ�CQz)�A���3�
��N�Q�
�nvJS�br���8pԆD=L�^2�k��V�S3��3��`Yߣ\E�8�!L%����q(�T�漈I�4 n�-��&!��a	}a��,��� ���Plu��O(�����$r�9C��Iċ=�S�*͑lE�7��T�M�ڀ~� P߯�Z�PN�7bQ�~a�8��"�K�D�_�i���Q����L��wrh (�mV��"��w&�y�X�<�u&so���}��z��C��f���g�"�!��v�/t|�G�lˀ���	�)��Ӗ�Y���oܭ1���ݽ��0#��'�'��$G����yk��P�T�k/X\�(29�j4:���sI�d�y�^w���ݠ�)r�
H֊��E e_l�t�<��x?�PWB��J����^H�F�dQ�"S=r�Y*�����~N�Tx�?B�A]Q�[�t�V��:DKƛD�ϟ
>��|A̩ �X�:�Qۓ�9Y�9��������2�Or�	ь��[v?�6FH?�b������-j} ��o_��R
s3TTV���P�(iP ��\��4&���mY����㮫�͉�[�`�2���{g֦.�m�	�ј	�!�tPc�Ј%X�t�_�!ԞU 5+@ݍ���j�NI<t��,,f>}��� �/B�U�%��4��H���+<�sqzN{�Vh��]�蓽|��z�t��ZWO,E���X���ij%M�l�vDӺ�.�߼8���a�4���ںoAl(���X&�ΎU�W8W�B`H��f��n-���֟�JuX9E�M�����֌����R����%#K��UHG	0���*yGY�l�$&���jSޟ��G�7���(R*X�!X��x��rX���w��� ��|y)$J�>!Z9�ڐ���s3�$��T�22��Z�6�>'R�R͡0��v��p��* 	pe	V�	��M\����|����ǎ�Y=���a�
^����3�� ����+GW��z�t����s`%�1M�i�*o`���I!	8]AR,n�ג�8WO�+��2h�JD����o	��&�7<�i��Έz�tC3\|n�5�i��xv<?Y��D�QD>��kƦUp��	M_��@���:�b�(���	u$�#Y��z�B<�1�� V\��u���{z��{�.(�� r	�F��9���)_b[�C]?1��g���~���2��47��˿��nH8��������T��{)T�"A߼'��VK[�1�_
��e�@+��}��.��DT��x�Hz�W�L*��c�ߑ��|��4sG�/-���8ܦ�q��F��p�ZfM#T6%ڸ�s�i:#��!�	 �cs����}DJ�Iy�Y�*��h����+R��أ�mJ�$�*0��ɵj^
�K{��	����Cj����p9F��
E�����3������_*�\�ȩ.-���y^�-�K�����ȴ<�BU���Q�b����i�=K�wԺe85%�90Q3��2���t_E�t�����-�,�Sc�(H8���'.H4E��)�j�n�v��#V'��N��2˾]��ĉ�tP�@�6m�P <h�S��X*�6�����;'jE��8�;���ط�`�O��j��ӏ��j�dy�>9���ؼF�6�m�� �>'��:l��nVk��9�g�� ��UP���9Z2�E�zS��3^�K6t{\�@I����{�d���,lin�䓕C���0�mc���}wB�(��P	����ZPJo�g�(���JU�f<��F��ڒn�	�4�kCv�i� �w�d�����%�4-0�E]L�#��X��5j�-�{9��e��7�1����J�pk��W]�k]��t����<?m���o_���%A�jW��c�k�p N�mc2D�[�<8�Qq�'�Q���0i�᛭���Yd��<�
i5s3 Vt
�6(���8�K��v��m~�?��u9�dU*a����F1��Mb�>�ս �-�oz�����+[��$1m2������_]-Ňk����c�R?�q�}o�3W���
L-
��\> �^�B`�o4w��Ϟ-�z�5����&l"R`Hܝ��s��K#<�a�8v����'ܒ)�|�d��&��[�7�s��&\� �j��ll�B	ãg#����I�UbE�8����T��N�=�G�Uc.ؘ�4\�mB��W�*gš�y�M���v�R�R�h#�i�%h�9�1G�N�2��!�F�fz7Ȩ� *o�b�d獑KN��C�f�1|��=�[f�ye]��ŉox��%j�~X.�L͠]�j��	0	�l��ס�Y��B�ęé@\s�O���I��<��>㭵m��<)y�n��eG̥P��X��Hg:��:�+��R��H�J���GN���HȻ��Jf[�#��8Kq�8��V��jW\�h�վġю�J"w�?��`jT�Ea2�mG��!Rx�\��~]g�����`vI���Cwz�o{��Ta�eڠfH��V�uiD�:.hh��(k����$���oTq�шd��I�}t~����Nqn�J��X�����J7����4����Ob������DY��ֿ�3@��P=�j���T��#������������*� �)����RE�m�_�*��9�"��m4};�{3Mą���k,�����C�[�q�C�k�\�wQD���\��J��D��2��)q��fb$�92��j�	�$j7o�����s9�^�Īa�A6��J�e��pڎ5��+1��ZnGl��5���}�Wp��WN��$��?��{TD��Qa��/ �)$Y��/h��;0^�����X�����G�7��3&U6����`�[���7�n��?� ���A�6�'�Ө�����Ѽ����"C�9C���l�8 >�y�<��Wl"�ps���1��A�]@ӎ�DuSqS��?�l������A���c��S�(�*������D��MԀ�x^@ �K�p\����pc.��F�}��6��0�mj����I��q���,���{
_�!};Z�ML����J�w�[�SZ{V��#��p��yY���#��l-X5h�hbKq���7T�b��ǴR�2��M�vcqط͇r���� 	4�q:���E�����>�\N����u衈Bb����C�kbd�'�C���2�u"����C�M���lj�]���!�p0˔c�@�؁�<�8o��i�s7+]��	E���a։(��V3Nl�D�s��,ʋ���m���\f�+7���Ӵ��4b�fe���,ױI�檱�:�|��*��{� �K-ٹw�:Z�\H�=�X®�d�M��g+)���O�`n%���Fp'?k�v ��({�q�Z!�7�z\�P�Ռ&g�#����/D�ҷ���ě�៊`����\@MM�h^���)�x�?YQ�4�DN�&0�j`�v4u�1=� ���+�T��Ο\��^���	G�����7���HC������[���_G������H	1�Q ;x�~DB��Wl�ΆjF��ۭĳ�.��X��r��[b�q��H��F/�����%�9J�a\�*��ץ�w��*k���&����:T��	�h�s�O�	�e8$\/dy�؃��m���u,HGb�{\�)�'�3�Xy�X1Ck�Ä�6��^��Y6��֩?푳�ɲ�B��Mv��N�P1�k
�2ރb�h��"�>�3^���%c��M��;.����~F�#�	IӬ�S��1���M�32�n^�2�nk�_Rv������R`#�Bx۵D�LX1%j�'�}���3γ-�W��M�'���9��P\�aU�xOFS�-��}�k�^�)D��e��'�զ7'PDD��	�\�Xxw���,7��u�?��Bdq��q����;����"�7��<c�o�q��H�OU��u�W�iWz��`�(�)>���r��E�c�趚�j��Ɇ����0��&�,U犝my�p�.��p�N���x��ͫ�\jCݑ&�?y宼��G�ǁ��I�� :\�s�͚��Sca";ǆaM�l>�M�����8�c$ɗ6`�-á�%�{�[Ս�����4�SnF��:L2��3�,���i��|N������#�ņ��~�%�z+���C��}�;J�
�8ֱ`6�p��NS����&��M���ǹ������∎�Ŕ)e}���X� i���H�ȣ�1�jّ��x�� } ���]d]8\��T�DDgљ־:4��x��)�Z�gyo}������;��L�cHS���"�+e�����XQ����z5���4�n"�-�gڱ�/��Y�'*��)��)$��P��!8DG��5�`!Ho�D���㴣�g1��U)�����ak{Ô_�b�Np�F?�"��b���\j��
�`/����^��t0�1@6�Bx�����o����d*��\�Af�%[�Б ��r���C~h���V?!,�Y5W�2��4z��'F��è���r��Q�9����vN�(��E�#"Z[�nne�@H&���I<��`��1u^Ui�^�y?@GJ�2� b���Ǥ"���%������Y*�f�׃�����{��z�J�ki��#r�z+L%!Y�l 	˔x����MCa�-1�#mUʦU#&l�鷏gOZF�O�Xe�N� �$(k�b�-�Ra���'�>�.�V%8r7+�iU'`xՐ*q)5o�w2��+�?/�ˈ����:��$ 8��e[O+K�4�=7�pd�PE:3nZ��ȩ���~R��|�7R''��s]NyR2����V������OW~g��/S��������l������8L\��Gc�ET�0�猟OATDv,v�p��F�΁rd뤳^(���>OI85u��R��$g�!�4k�i,0�G�Sd����M(�=Z" D؍���D��3o�x8�k�&)6
j�$#�$P�&���H�0�Nl��K�1����C�ɐ��(�t���)DK��+���@a`���1y���o���:i�F>��:��A�+�eU3�"����O�G�4�`�'Z{��y�Ҁ��/��]N@.HS��������j̡�P���r!\�eꪓ��@49�jm��]&)�[XA���J)��B�Jg�;�.8��u��Z��̓ʂ�����"���i��FfS�x��.�4H�7j�/�?<�?�7�}ң�k�R��Kiȫ]#��G'��i}"�z��=#[>i����
�����TeD�ݬy�8dȭ���B0l
α8�Ͱ�9F?�2�HQ����"j�C��uk&�	���$��u�#-	�I�T��=ꏂU���3����Ү�2�Q�,���tv��6��i}��p�%q_g��5��ʸ��F�7��=�69h���5�Ԯ|�w!��$�"��X;37N��p���W�����E�cO���{���/�#�<b��k4�	�{D�NL�Nʓ��q�R胻p}{�T������K��w�<4�����x��_�ס�4'D������64��VP���R���<�UӔm��u�F�Ɉ<e�s�W����L<?E(����˘���	=`!�.=i<�eUc���s�{fw���z�B�ٳ^l���Ⱦ�?�~����Y�F��6U�3e��[h�A��vf�(��T�-�Ldת��]��]�6]���g�1�A�)6i�f��џ��V&ge>z�K.�� �N� ��Gp��:�x�ru�����Sˬ���D��;���/
�At�|�#1'j榑:D��-���j��ϒP����̈́�̯���6%�~n���9��-���)��w�fq��a%%����$���mt�)'o.#��|7��id���S �������{��O�z6��g� �cBl��xv;M�nc�z�U�!��!�k4�P^)�J�,��'L�	�7�QW���޾�/�]�U`w֜�4��}Y�<tp��L�o��-BW���+\>3�G:��6
V	�~'�[]���1-����>�z����m:���p��Q��E��	��&�F�+2�����	������ufu��?�~�q��v,�������H_+h�B�\#�0l�a��r�����U�X�9��f-� ǆ��^X��;)u
̍�a�.��|b��#��� �W�K-f��L���~1��CҾ������$ހ��k�H��;�B���p��?y�"�m!��Ej4�\�߳%t�c�B���*k���'�1���v��n�����y[w�ҞwO�u�����>��j���g�
@c���_���[8V�������ߩS|z/�[ú��#�="�2²+���S�=t�D�����\�>]f�]�OsY��vE��g���8�F�����5��+/M�U��|TAM	�d���S��@f'�|�"��);�t��Oዚ��/[>tɷ}�_ITZ�Ii^Xk��c�yd+��ct(X�j��T���	� �'�����J���o�]N?��B�ӾYԪxe���~�},}���*��[+��A�}Il����Q�^�0 �į�:0�����y��~%[1��}C$��f{a�2l��f����d� y�r��#X
Y��h�Z3~8@�� �^�v���X�j�*���:��4ABZVd��� � ��?�n�̅G�ɇi�EK]�{��RN_Tf�ů�����Iܳ����t:i~������tO5>G�
��յْ5Yة�;�:1c%9������=�PH�m8�����+�G�R��
�8�l�c`�{�A4ȼ'R�|�:Ygs�-�����e�/b��߭����Mj��Z��9��|+q���/Fp/%��%H�m;�P� ��	�=�&@�H�!�x�W���ʯ�"�����1���.�55�.)�K����;�Jɀ���t]���O/�e�8՘}w�!�>�Vr��R�pD�7&�����&b�&�raY��E�āۜ�s�&�N��`��KK;n�Ё�h�3L:����b;�1v��+����.nі/��\�b��Y�i�г>$�Ը�����2+���F�h�R*h������ȥ�F{��zm����N()6f���'ர�<�¢���#iF��@����A���_�&2�����:��^�w�W��*�����?���(�g���]���,'Z�u���y���ʬ�BT���0�0BI��J�'9����c�t��WV\�2��@�^f�T�}^��P��j���T������u�SmPfñ���L��C?_��]zJ�� ?D����;�M�;o$�z����Uk����tB�������
+��?�F`^E�$J�W�]4m�D��Aa��D�D�U�/+
�h�� �l�u�R.SĖ�=�@��7���T�-���}� �Q�!]P��q6��A�T)X�B�5ӕ��6��5X;����2���9xչ"-���r;��xcɅ�gI�"�����~��n[*d��-]U�a]\�c�_v��p�����Q�U�#��HI�J\�O�ڰ����q���p����>5������i��#�o":p�<3n�)�taXz������ޫV��j����dL� �y�^J��Q,��l�l�)���?�����/�mgH�3����n���&t�AO����,IAc��P�3������N����GB���R=�)��_�H��^��m�:��
��?�^0ԬФ��ң�w�YH��gn͓��Y���s)CN#y)�^1��T}/�9w�R�!��"���P���d�=)�ZA!Ł���c���ܳ�9���Γ��7�ŴH�Ȅ���U̸�3�Ғ��cA,�"tރ���
�������>��C+ŏ�����a=
N	P��:���ٓܰ����o4����iY���r۬;��)��C�xS
��.�Y���y��Q��ڷ��%����ń��"�R�F�Ĳ���v6MB8G��!:hj���
��W� ��|�W��k2���� ��r,Tiy,w�#s�&�q�+��xGI|��d�^�l?J���b}|�pn�b�6�ؕ}��aY,"ƪ�먧�FÐoha�-�m�:h��V�l��H�$�$�K�2^P�mNД2�H�m��Cj��P�����@r㷄I8��˞�����F�^��1���$�9����3���){�B��j�C�0 pդ�/�Շ��E�A~�HY�Dɲ m�m
o��6�"7aX���^����� gV���7Q�H�1�HH���Y��41��_��ܸXV��
)���ѐxڕ�	�>CUY�ʒ��C?ko7��ʺ�cQ3��T�P�"%lM������Ch�c�$�Rl��M��uu�} �Yh#drpL���۩ᕑ⢺D�3�>�>��	7� F;!�Id�YĖ�0E�a�&,���
��u��H0�{D�G��S �m��=�N��� ��w��C�t��w���:E��1�Gܷ�����8�W�:a؀��8meg��;��]�h���^��7�S�n�l �f�M��^����Ю-��'s���3̞���OG��S�d��(q�G�c=l�9+�8�����ml�	�/I�VM73���ɞ�b��P��ѹm�����Y��Bf�E�����]��5zh�|���[�7(L��#;Nx
�k�����G���~�~GlmϝtS�N �d�+��z}�j�6o�o*$1R�=]�.L�K����$�@��F�%�O����yj�����(�,^E�#�w�$Y����G��j��2�\\����-Q�m6㓽�vl�nY6����R���Ep**��b/,(R�>J����֌�4�`�J�-B0��ZV�9��njx��5l��� �
7�'nU��<1U�WʒGJ;w�XHt�̈́ |�ɱ�ϛ�e�_�M�n􎦥�ͿG$�e_�[�#2;Sv���\���<�"*ǔ���Wh���BFɼ���%zi�z��@@�V��@�f�cOP�����`w��b���4��X$�5�}Nk�����K���M��F=�[̶]A�z����mt��w}�����&#�B��f�1�f���AnB00�n�3��ë�?Tn��R�G�����x�mE�� ��ءj�����A@~Ѩ;o�4���Y��.��̡#�mP.ϪjE��j�ȱ�4��F��̞��2KnS1�����?�Y��~�eY�}1�V���	hv��鉈��9yd�"��B�i>���^��g�7{�/�b�p��&��
@�l��6�~�,��~~h"M�������22GCj��Pe�H�__-����ֳ�W�хN�u��P0<Q�v���p~���I�[�������=+�V3�0�A8�T���~�(&B�d����u��("E��mW�ĳ�?\�˽4?`O���ӱ�i�y���F�`��I�[��cږ�qF�'ȇi�՗���z�9�@�Z�9�j�	�E.��a�^�k�L9)�d��M��P�=�Lչ�:�r�x+�*���p�z��G�qjȰ��{�Hq�s���o�z��~�f�q�n�ڹ�E6�5et*�I9���[:�孌0sC;�~�˿rȅ��!m�~ux��3cL��ǐOt�g����#���C�9��΍+1{#l�?
�9L�,w��n��v0� au�3;���T�V�������"�L�H���'{M����n٣���
��O��i�~hl+�XR���)�W�j|d�֑mw$�GV�2듿Q�]�` �.������X��� *���݅�FZ{w���j�IB����q�Pլ:�v;z�7|C����"�P�����uh���B���c'�FU#�A�k��ul@���>���gz��k�^��F��3��txЪjA&�c�����j���7�Eq~�*�1 �?�K��N����<�["������`�%��}��i��-)<t���X*�1�4��	HS����4�W��E�|yGFc�!���j�hYǃ��V����α��K��y=�@n0@�8�Ŋ`��
id3<�t���FvXlz���B�{��e[���4}O��h��~A>Tή
@E���f��q,s5�Я���/�4���Yl�R� S1qP*�����UY�(G��;8�yU)c�*�9M�R�QBS�����Yn-k����۲��=��S��|�}#�X�s�5֯����T�~^'?Q,M[�%xK%>�b��yHΈ��p�_���d�����M���J=ُ~<�-Iz�REG��������f2����ym�K|�4 ��x#�c��h���-9|rp�����a��=�{���B���	d�Q>�^��U������A�ʡp1��L���/fQ��\Z�B�#�]�X彟am�w�ٶ���\�7wg�.J?✫�q���ͶC�Z�}a��y�ˌ3�m]�)�#h�yl�>�G>�(p���c�6����ũ�v��o�%koz�w������U�^y?�0�eq+���7S�Ȓ%�G�i癹_��R��
����ۡ苡ˁ���]�%����}nK�������i��]�[!s��������;b��WA�̌��4��훞M�7;��#m� �
ɉ����`�� �LR%�	� ��*ء�+�OT���p��	�/v|9�w�"���ң�,��X�B�39%F�yw{}0�nuBqBHC�@�=�~��;��\E'�FU��|�gg�Y��
|�����L��݂TX�Ĥ��Į���?ڊ:
r��Ƅ^��8��NCͱ�]h<h>3S�D��	����>r�з����j�Np�eu(�!)�B�đÜ���������̿7�E����(�S��/Y"�V��"���'%c�	��Q�<9-&x9�G�Tz��4 J h�Ԓl&m^R�F4���uK!
����FϘ��a"$Q>,�lǼd��f���^��u�/�럧����ʞQ�=���I����׶�����|�L!(i���xF$����>�o4! �6$s�^�O���������e���ӆ���>�����k�����T S��N���q�LoN�M����;� .g�KF�����U��)�Ñ{.�񭧙u@�����~C��ۄ�u�L��@Fj�)�L��gJ�y����`�#xW4����q��~ f+��e�e^$r�B~�&�s��Z2�Z~�
��&6Z��Kmc��jz�{h#&��r'�ĘǾ�yS�ܘl���9d�
;L��E5'��!8�f̬U5ଦ6n-�7y���ѤȤ4��`�Fe�2�C�:�U�y�'�d����aYtjU:'a�bp$8�I6�l\�c�[���i�����_��I]�be�~����ZnG�^��Մ��Γ3�W���ަ��K���	VDFMϊu3[��r�R��uY����[C��� ^��36H���s���c��.�I�}&�5�QM\ D�E)��jY���l3$�-�j�:�����$���V �0P��P�/Ӕ2�2ս%|�b5�.oV>_?)��>�!�w��qKo���P����0|}�W1��a-W��U�8E|zp��P�[��<5��ku^�Y�m�K��f+TS8���cT:�4���;K)��/J���hS�\R��~7���9�P�]�l�;����l!�C*��64�|j;�%�ST>�;a6Fק�?��h�0����HG'��wj�1�gu�m�#Ehw�ǆ�{����X����9õ�X�'�e�7��<t����kZ�dኃ�!6 +
����ɐ�ZxM�7�����s��X��z�uw09
�V��$�u���ˢC��^w�9�ְ`��ogB� ��u�?~�-�iOg�`u�M�[�w���VO�\�%e�>ɾ��=� 
+kO_ S
��Փ����Y�SAZ�M@��l��}���G��Yk=䍂��W�����.Oٜz^"���0q?D֔`˃7���9��ϳ/L�)B��)t�`������-9��'0�.R�>���BWv�q4�i����z�zkNϦ�K-���0�-��	e&6s$��?r���(z�?ѥ셲�H�	�0��~�vĩ}���7�um��K���4��W.b�����J_㤔�G��V6�ݶ�LȌ��e��L�y-�t�p�c���uV���1��"��{���2ټo�U+��O�P��S"ː�G%\��Q���s~ZF�����!�{��8/�"�W+rV�
�e�X$ۅle��-@��ec�U_�$H?B{U�s�5(����W�������{^'fH=��iDZ�(x�c�% w��֘�Ώ�k��J���a�>6�~�6y�=��)):/I)�b��Ai	;}sD�7G�����:�[4�g!;[i!�ZаD�e �"�����&�Ӯ�N�!μV7��ߍ����Gh/#[��v�#:�h��F�3��&��w~zt��Ki�3(g��,+5�Xګ��M7���9~eIO<n-jl�vϋ/���dWϺ�P��Y���W{��Ǟ����$C������K�hGQ�PN�<D�̰_�J4���WxfX��PF�� \Y�\�
*5kT��ō�o������颊�;�fG��nU�/��t�dT��Ĩ�6E徎�ۻ9h�)��J?/t$��p4��?�5���7�&�PǌI�ɽ�����q:�Áed)��k�41�B%���q��2`��3us�A-��"_���	[ӂ���	���ŏs�w��\G%5�( Ӻs�t[q�U�4k��l��Sd����FK�1�S��R�J1���~RE�(��!Y��M����}�ܤe|�����P������t~:R��o`Jo�×ն:�Ť��xM�UΓׁ�x'��� Ϫk��a�_�� �o	�����qi��Ey�nf�3gz!SL�ӹ*,>z퐍��u ����Uµ%\}·��U�se�ƹ�7`ȹ��;t^����s.-��B,��e/a����{g��Q	�w!5� �N�"ٚ��jŷ3!�ö���ڣ�^��Y����N:/O�E<i!�ZMQh��̏V�mE��}��Wmk�n��a���l��HI��|dsm����>˥&A}QNiX�'�x>E�K�Eed��T(�K�݈�����_.���=����;UԄض�a2�rZ�h��������&l�>YϹ$��ѻǴZ46�>���yl�ؒ'�hn�>9� ��V�������S>$r�����l7��'Ȇý��}I�, �$Q	V�S��{�aϴ�JZ���hR�
�c$��f�ⳋ��k.`���ʈ��
7J�,A4 �Z.s�nW|��R� j���p�'��S�x�n�)��g껍�'Fg� �V��E�B���	LM�t~���4���]q�l�{?��[	27���-Q����Ԟ.o�I�q�}�v����u�0�?f,�q��-�`+q<�MuM:LAᣱ�9�%5��3>΢ڇ'�o�2��4�d-�(&p���H5ԕ�g�d]&,?���@0h/:�P8 ��T<-�_w9v��oI#����{�mw�fkOu�C�!$�Д�z�J�����}H���?��4o���.I`��a���;x������w���u�����`��c�`��������������	v�q�f]�@��kG�{y����
��S����.�
���M��.<x��)<���K���Qu���c��i�Q��a1�Q�]!���1 YTn�#|���+Fj���-��"�1��"��|`����`�ZŶ}����:�|�V/%���k��}rZP���P�;
|�T"DC9K\
���|��!�EV�J�qZTC��|=7���!�EPF�2R��P=˗��In��J�^7M� i�-_�Ϻ#)]^p�R�C���>'1�#����&�Wf��5A���$)S>����$;M*�s�F���s��m�G6~�V�b̫�K­1B�T�u�>�e��0�f��Y�8�{��I��@�� �W($��`k�]5�!�Q]��� 7��q0�
�q��"A�����hRܼ��〟�ޮ�l�����3f��=� C�>�#Fu"�bo���8��rmY�v.���aB��` ��Z�'Ɉ������H����-���N�|ӯ阚�~тa�/e��
m�nT����ףY��>��#�A�^���x���<!�d�J�0����H�;}>�P�i9��A�&Τ
ݍ������zJ���aS�\p�!XNc�c�cʃnSi�]�B�ɢ���7��
r% ���p%��zVa^���{lz��X����&o�g�`��YKj���5��9bZ��(�ުn7K�u�1�*3��Cw<IB��GX'v%ؿ�q���c���)�;|���)<=LM�({2��-NT�I��B�l���$������)Jw;����������sh:�ix�,�q��t��1A���j�0�p�*��F�.�og�./���5�|�Z�KЩG-_���!y�c���X��o�bI��\�bd\u�A %���r�6�������p��7�H�B��o�&�4������c�+'f5�ra����+�����7>����H�$`�nr�J~���"��)v��
��IY&�s'E!���FT�*�Y��#�9�F����i)��_��m1�Q4Y���D�59�v��%�?���;&:I.8O�ic��Д}ی��(�]���F&�T��(!j�ª�/$A~3����������)�Iy���SHi(M��9���G�ͷN�x���7����*NQ�]qȘSZ�M��o��,/3RD�O\�ӻ��)lu��v��ԃ3#I�B����E>�1UzB���#��������b���b[�ۃ�Q��2,$
\H��t�7�3-�!<9�nɚ���Ӫ��65����n���wr;y�S��9_uGʌN�p37�*�He!B[�c]���Ǒ|L��4e�����j��*�:G�E��0>k������7�5��i;��C�"�A��ghp�W���)�z�-o�6����K����Rh����;]`���M����<Oc|S�PeL��\qI�g��X0��Oj2�g/���z�:^;�����߻���֝�&�܀������O��&h�(%���?�[8�e���po;�;�<ǈ�ţɦW����0I��-9fI���i�#������y�hٕ��4�k��%����V��Y�'�����T3�D�vBղ��2�mܸ�����y�	�M���|=B���tW�A%$	}#T�W���Y�ŨN����	�Y�-�M;��lfh0����uW���6�qbW\.F�̆Q�Zbg4VT�q��j�Mk44U�k2�W71̺?�� �`?��~FN_ˎM߳����m���\�����"��c0^7xp��x3�n��;>��I�\��ߪP/+8��a�7����~8���鴗�S�*��F�_d�Ӫ�/�Ϫ�mI��N����K�K��'���T��N��W��o�%�%��ջT�A��2H؜�9X9m}[_k��A&�L�f¤�i�̏G�2�9���z�{�26��\�vI�7*1���v#�Se	��q���\%3b�r��� H����Z��y�n�����`<n��g-
;�^s���1�4��q@ƒ�/������H6b,4��޴=�M ��{ ����Q���N0+�B۷�f�`��;I�o%�*�%�������>G7�D! �$�5�qQQ9�HN�zz���
O��(�G��=��4EL�FQ�*g乃s�B#*�H���� �F���4��T�M��	� &^�	l���թ�]k�U���{�x�L.�@��ДU'Y"?��ň9�Ub�:��t���j�lj� �������n�>�u!�.q�Z����K$�p6d}��0���JG�4�ِ�^��l6Ll.�(��n�2���Г+��<s�/�T�>�q�.��a�)2n*g�4<�'0��E儸Tܜ<.x���]�֌?Y�8��M��x���}�i)NAA#��Vqb��/A_u��a\#�퓊����� 
,�(��K�_�!+��^�Ǉ�\t4,>����$�m��Q*4�z��#��b�����)���3�!}'r�AypL(��rq�7���G���A�J"�\Ut�o~���#�����Bj�pV�d�yT��IA���]�8�	�T�<���k�Owh��,��'���9�N������k�
FH��!��'���WeV�D-�C# ]@󲢒Ma�D�cG����ސ��%�
z5]�W�$$3ÁQv�[.*^,#ղ���kN��:��~PJ}�g$j��!N��F_jWE/��N�F�i�\���g�u�*�SZ�cҼ%�n���mc���C0c�o"_�EBB�Jp��A��N��fK��
��5�--l*`o����X��|�B3/� �Y
�!ra`�J�.����h攞i���e��P�{���Ր#��RKy�k�7`�SVs~��퀽����Ucd���0~�Y��G�.XA��O���,�w����E"�J���t/a�AK� �s��y�4��i�Zt���>�ki��"w�w�D��3[B^veJ4pgi����2�n-Nc�U����h����0[�Y�����]RL�gD{Em{�%�i�Dל���3{G�ij�4Śd�	U;���5�Q��\�$RDC��:�bf�W�&e|���<�M�v�7�R��~2-�y��� �����N���QUk կ�G��Xˤ2R�#S�;�(�g�O����!�?�9�M�(��ͧ��8�!�C���-�xx���~!)�(Bf[�/7���[�KR������Ȗ��޾ �Q���Q�&�.���$WmF,�����S��Zl뛨���M��ꈴD�����:kCH[�L²ټ43G����u%=���KA�Ybl7��#O3�_�b�P�\��1� �ԅ��E�����9�?��'�an�6$�B_C��Wf6�=��3�i]�I��-|ʷ���Sw���_ &Р�E�g�w6H�H��ԩ^�v����f����+=���N��Jaζa�\�1�&�57���Pڙ��ޏ�{I������7e���-���YRgt��)��B�Uǣ|�x�Z��ҳk=oA=��w=�A�[GA��u�U�sшzn�%���~��4:�)\X�>�B��TM�a$2��2�f���%�V��(��Z��
�#��ͲC�Ul��Na�"�����I�	�23��ɉ���X�ʟ�$*r_?��\�B�#�Y6���ӳ8��6*���p�!ϻG��X�Ȇ��E�En[������tC��d9^�O�c�H�ޮiQ%�٪��%��I�%���F�wn^QOMx���o�H"�p�3��-麴��ij)��I>j0 @�6,�4g�(�a�X�j����$�Mt�"�����S�ֽ���^��b����+����n����Z39?��R5em}�M�� +pB\�06�~�Zl��U�0�Э��/x�qx>:�jK���o9��}^� ���"%��ʅ�L�@ż�_�*�!m�
�4j킔9��Y��O�U���ΐ�p2}�w΂AP"�k�@0�Ơ٪�S�&J~���
��A�M��A�3���Bsl���#Y����ʋ���rs?]�zlr����؞R5�� ��n�H��6����5�Wtf��k'�M��˼�Ky��'�Č2d�"������A�����mTP�f�tѬ0�ԝb��E쬋�ɛx��鴛E��u�fr��Asf����)�=+eM��z��C���Ht$�^�N���ƾ�|�����^�ʤq/�\k}F�e-gW�!�42�Y�JݎZh�d�(C�o�3�o6%.tT���H��A�X��!|����p���:Vc@�y��5*�+JidL�"�u�������*T�X5��	�,|���kۭNY=�
��e�CW,�����8��gx�pٹ#%_�7%_��1w���Fn�&�X���=���jߴ���5 �s%Q�
	��,A�i*��u (�i�Zf�=l���M�-g�Nh��@X���n����al����Ň�K(��]XN=��e����:���Snw�B�5+���UA̟���;������vg;z��I�,2�9���k����)�B�?�^��P��$�I�_I������m�$�0�)��A4����D3O�;��:ZL fv���v�@u�x��t!{1U����cQ�X%�r�|M��z��f�:m?�vB�lIܟ��T^�2KK��R��opui�.�_8"�F�-U��0�U}~<Z��l���Z��C�/���D��s�Je?�Zv��Z�6
�4����ttE!RbDl����`.��E��x:r
Vb��%R�!Ϡ�'�%��C���ݓ�a��v�@����M��Gnh��1�V���:�����]�h�7[6�'�{�#5�OGS�U����s��h������H��v��{����Bf��iY��&u۲?�h�0��#�M� r<7��N�֚%�ņ��VE�T���m������Xx��k+�X~,����@�\�0�ٜ��
��ׇE1�q����r,���w�z�qq�&�5ntc�\��MMP��Ye��a�V������IHV�0�[ZHkj�y	Il:�몾��"��j�m��l�'RŸ�v��}�*Z�[�
��C��@|��܎`���ٌۻ֗2H����ꎴ�0���뎪���xݘ�r!aD�Ky�7�G�k��j�� &��`i5_Y������[.�ʃ�4��� c���+}���E< §8��ٽ5nN]t�4�q'y���ۥ���.D���6��.6hЌ'M�b*�C���U�� S3GM��spW����OUN���s����@0��ӵ�f���{�>^��q|e�����!��\�L�:�ʘq��$f�']�/�B:�*����/�$�ȡ�v;��(��2cDm8*bB��aj�H��4k;�..
}x�Ab��J\ѳ�g4����%~��T+T�����ڷK�@v2�p��AZ:��5sԹq�8�&��^�d���*��Pd��/�h�F�iy�j�{Px�~�}j���Ƭ���cEA�D�g!�F$iK��J�wt"Q�V��<�N��J=E�8w��xԎ�)eU��r���"aZ���U���)�;���e7���Z#i8-z��_��}�Pe:V�,1��2�B�'M��;��('K�m	O��C�0q�x�'�ߓ۟�D(e����Z���*��'�c�h�{�=!�G���V�A.�2���Cq	|��z����ZZ"xπVp45�B�"��J{�Rm�������sF�����3\Se���\�'�4����A�I-��ow^5���ھ�mj��ڬ��^3#Rl���������ǖ����Ê����_g�u!���}����sR�F�!:�����a��r�<�ɽ�����'81�Z{�Ɠ�ɺ��xf���@R@JP|n��� *Z�ڋPN��I�:B��� r���h'��������y��V$D1g�t�=�'e���Eb�S��p�V�h���FnP��sq�U�@�Q+�(��������p*S �#�ح���#�/�7��]$�&|A�Bz	��R(L
~�^�9_��뽾�/����n���'mk���=��jӬ�E��w�D�Zz�����h��Li��ߕ���;��5��t�X� �tP�A!'�4?�}v�HDL�f�	{�����$-vv؟�xو��z���%���	���ؿ�V������jI�*�:o����T��8*U}�m���?0#�����p�-� ��Ðf͆AC�P��x;h�-b8��f�G|���L
�ն����	�ɸ5�Q�{��YI���zQ�NTl
Hw`�vY�1��O%�̸�F>U��D�/B��m"�(a&ÌWԤrxe��%�W��!��\}|Y����Jy��}
�ot�l}Nr�B�˘����p���;��W&.g��%pK��`��/�tg0j4{U5�I��W)}�h|si�Q_,��om�u*����ƺ��#t�O>9m-�OH>���ۑ�c!�wW_��I������&�U�9铉�TA�>��j{J�xF�a�7���X&I����-@t��9E�~��U��d��N�dŢ|"�>���J�Z�W6R#��A�C![����!|�C��"��L��[�6�y����U;'�,?�.�}���O�.�kX��`���3]i�6���*þ'"�s������7Y؝��YU� 	�M{���hwܗ198Ht�ǿ=�;R |l�6U�ƚiҏ�j��!���	DCx(T�9N���jf9�i!ˍ�cY���@UG���|t�s���&��?̋����!=�tE��Y4:�z�|T���$�.������lB�V�����\_�v)f7�dU��+�KR��z0��7��cc� �������{bx��~MTS_�ڥ�Ju%���:�{��&W�V�{���0m'����h�u� {w�1h=�D�H����<�wkM���Z���z)���L5�U��=z�|T 8�ە�Y[��p�"Ý�F���{���J���1H:i�ץ<ߵ��_�����ӯ�T1>�g�+��<)�1Wݎ/��*/���͘D�9�	���9��,s����U��ͳ��=.�i�K�$�-�0cVF���Vy4-j�l��l
=����̃1��l�i���L3����I�� ����䄊�Q��9�x����+�2�,�<"c�(\\�:.��S.�{��[ü�wg��7j׉�	�'p���k��m������W�1�����چ/ӂ/�źu��� q�ZTY�9>j'R����.=�PnO6A���K	M6z`:U^ݕ!�0�aZ/�o�>Ĩ�	����9�1D���p	Q�9�ظ-B4��Ed�n��T�x<�-`��@�|��P��DM?C��S�'X;�٣;݇��C��h��S��!��:��3�Yì3X��6 "{Nu�����?��_Mtw��ɪ�3�1����풜��[`+˘
l��P?Ҟ2�Xk�Q@�}�	�~騵���x�� �8~�o�y�?�ϣ��-�ţ���@|�yƗ����z���j�b�(鳇��P��&d��� a���,�HCy�t�GS)۪�Y�r��א;���0Z�jf%���!
���$���}R�z�fšPX6�0�s(Ba��j��N�|Ĩ�n��+�\� �ȕ!wT���s�
����c����|��&�T��^J�0�l^8x�n����t��jpÜj���d��Ӌ�'�9���]oG:��닢���מ�B}�Y��d���=Q�L�����s!q,��?��/�d�OLntM�!m�U>ȏ}	�0q��ӯ'����0ѫ�d��Wޘ�?L��C�ɡ�2��8�G��Ut~��Ta�����3�r��尻k7V��09 �'�0-t�'��6��&�9�Q�sF�S�g�'2��
���^IO#"�"�R��:�{P�����#u��	D3���3/�,���XtD%��V������E�`��6��u�iP�i�����v�d29յaX�������y��1zfk�{Ρ�%�� ;���_�R��5+��	�2b��t�8�U�c��ҹY� 
�(�N$~���J��~�W���Zg�;k@�ղ6W�A�����_C�I�^[�r��m=��ǥ�U�z���dm��!_���T�b�2&j�!�d)��W9�*������s%�r�`�a-� 5�пj��"=�i)��Q~�9�j �"��'��x��"���!t�>�,�V�3O%o]�)t�J��ځ�M�5��U��3S�x�-.�-��CE�?W탷x/��9U��T����V��+����`�n�� >1�����`���_c��tǛ@r���ᷞ� 81�Q�̧y=�s��vz^�gpˍ���N���g�ǂ8G�b0�A�Me�8$���w�_��j(R��!����2/e�"�����<C��b%��B�Dp�
�mY}3(
����}l������>j�o��u�dDkk�<.��>��(�_J�R��6�:O�sw�&赮n����-j�Q<��c(p�fQ�F.Fp��j��R�2�j��u0�:�O�l�٨'#�KP��yu�pRO�t۴� ���rj*+Gw����0:���xʹ�z}�.�ٖ�|ŏt����)]�5CN\x�Lͤ�����K�.zEkK($��3?�4{ʉw��[�SM������'�
v� ?�v�Nq��mgc*����{Y(�&[�x������
�뢲�d���͛�z6�=-|�)+2`;��t��H��M��^��L[�P�uK����3��b�&wr�d8�ZC.R�S$�ݲ�3%�2�hk�8�R���
�Ѡ��Q��Z���u�Aמ��*�b���n���`���@'s����c�C4�����7�k�����jЪ0���JwSj�gW	.0{�T��v���I��J^�(�M�g)0�z%�{7-�=8��6������1�X?�����6�#2^��E�����ʝ�#B�дK�*����yyz��RJ��޽/�6��H���J	� m�H^yy�.�27A��X�����G#z����p1P����i�jC��;����(L��� �Qߘ�=2�o������5�y���mTt�n����}z���Xt���Vǀ���L�i��>p/Z��K,�Ҳ�A�u{�y����I��Y�?V47A'`lכGi�i'0 h��u�r<�9��l��6�O���Y�[h�s߸��#��d�h	��,�ݾX��CA:4�j��r�g��4v�gZ�lmT�ȗ���mR7l1�"��b�:9b��ԓ�=�K�e潅��l�H�WFy�L��w�j�����q{b ķx17�s��Zo���L����4�z�>'��j�
-_.lǙ�Zi�.�<HiR�Q��W��0#���� X���=Ҳ�eJ��Cy0㒶�.bϛQ�=�ܒɵ]ў�5 �ۣ�QmV����\_�n/��紧��Ix�'�T��]�Ƭ]B�-������fЁ��o𺮒�$|p��!��Ɩ7���T:�j�Y���B*��b��7[��C{=�^���K%9�@�?�ڀ6|)�ى
=&"~4���[���LH��Ԙ��7�Б4�}θQw31�c��Y�b��mBb�ٟ<,X_6��l A��p� ���n<��W�e�hQ�i���.'*QnQԀ��bW��`,rK=DǇNH��@��.��OrG����E�UBަbv;���Ϙ�����?.l��o�vL-o"�8Ɲ�����ZB\~���\��,�������2�+��f���q��p�T>�N=֐b���a�����he3Z=�Gi��8�9��z&�t����Y����1�X��F��!*�B�6ćf�*
���L��{�9ZdC����X�F�Hc�jA�J�,(�66����;��W�}��]��M���T��ښ�ل쯴x�3@����b����@l{�\i}�To@���{��m��{��O	�\�ҫ�'?�˻�k��� Qf.�mㄵiN��h��V���= �D�d� ٝ\��Ql�\��KS��`�r��Ok�(��?�q�������)��[�C��*�]�A�� Ԛ�UǁM= '�c�0�Y����5p9�E�а�!Š1B��Ƴ��nY�Ӈ03������*z�/v@�����Ll�Ywpn�A����"��`jeE�#�k�I�K�[�D�4�!1>�Ę
b���0�����wv_��EO��d�?�i9��K7���$�`�6�7:��.�����7���X����U�"s�����ւ�q<A��	�3���d�FG�H�*�`٪�s��QM~A�W�.S�(�c�Ǹ`�Ք 2�8j��2�$T~�I�[P�v�:Y�a~���9���v
��( ��mRv��\��M!�4�u�k�8��r�w��Wy6-DMw��g201�DŢ���'C��x��9-|�v/��Oa�L	��5���{?6�힟XI��/�������t%�/�ܟ}\Pǋj�4ks4.T��F.����~�@~��#��ibR��(�n�j�tx!�F1<�u��i8[�Tw��xu
!�64,�rAeu���� Ѝ�����O1��F��(S��&��	Y�QzJ�viq6z�Ke:�x�һc�������Zɒ6� �9G�8�4!�Pwa\� w��i<>F�v����=�9&�S�'����~止�v|B���d�5H ����1ΔKVn�����!���].���4�.)�!���Tr�M��*_��!	�EWrQ�m�!QCCkbn}7��ʪ3S�g����<o��18uI��\��5;E-�U;Ѩ�H#�48^\K']!@��N�W�a]�<1=	�*R'es���g�U錋T��t�
��K�.*��dNC��󟓠ˁ�~�#y�R���8$e���=/�3lÞ�F'�zD��t�aA*ZI\V�9�q�G)��1�X�Ii�h_1�!f{����'@�,�6�Im����/�����X��sJ]-�����j���G�',��ªM�V&�v���T�T4\e��:�>��5o�${�@< ��np�W��[T߾L�/����Y��}�e����E��?����c����������3�n=�ʫ�(/�s��3x�5cn��JPV͓Y���P�$��f��Ñ�o0�<�f����A�u�@X� o���C]9i���C҉��h�D�*���޳JL+��G���BF��zC��/Fb����Kd���ń��n��'����`�JJ��7�r0N{=$rҷ�kg@t�X�P�@�"r��W:)�ﶪ?}Cu}Z����Gc�S�ٽ$�f�i�Ss%B�8��"]*؏��&��=�䓉�S�j΁�����j��*^��n�.�|�����=xe=A�r�w�'*f�='��K5s���S4�#|m�ˈ`�VҬ�µxg���M��Y����!D;=ڜ�L�cp�h�|���Q��ꞵc_�X1�䆻>՚���uɺ)l�::D����i�'s<�丗��s��Jl��2G�� c�S��XAZ�0�m��n��f,j�4�z�L&�k�~
 a�8��`���S������0iQ�����q�f�$��
��z�9��:�-�Y$XU�������+���A��ͯV�,C���F-SC/�9���l������U�7������Ұ|�v�qz�;��ߒ�`&4=���@܉Q$��|=G��kP<F�r
k,��A���_^�-/��n�	�q�2��w�_�b�|���\<ij�o�=Ο;:d�k��^d���!���u����<�]����Q��q|�ݤ�څ������01�YΑ��Yp?h[c���!� �uȲ�s���pc�����S�S�I_��TM���o�>Rn���&���h�h������e7׭:�G���	~�i=~��c�+KC����
�t`��&2Lh=�ۿ$Ь�0������Jk5\yH�<�2�5�M�H�8�����1���ڤ����څc�[�u�Gv�Z3�=uUb��+�	�^�C��?X=Jj�#���yWN���t썄s�-��T�7��̼r(��	(��W /��:��(~e%Š�� �z���W�ƪ��ZP$��	�(����k�Qv0�p���T�le��i�%�v��<y�Z�� )��l1�Ul�	�zzR�[���Og�����h��9}V�*�ϟ��m�^�~��ܑ8�i��_��1!:�"<�hM��b���<-�?-4�ў�<S:�V+nۃQ�,%���4��4���e�O�'vP�S�sjb�R��-�[����|���	��܉xǋ�^�3ǂ����Q���*Pz�0?�/��A�[)�md�ࠏ~��نm�H�������=>Y��59kx���[Ke�i�ǜ�^�%���DSF���x*�j��Lf�S�җ��K�〫��jx窷�Ԓ�]��Z��Ӌ�w��׿���#�����UՆ�Q�����Ό:4!;�]�y=��&����"#�
vR�k�༭�����{O�\A�WAw��9v��,:=����Ta���ZƺA�P�e5�ks7�;��kF�^�z��h^�f�QX^�O��b��V� �{�x��DFɽ�ɓL�#���uI�º��:�)ￕ�:�r#�twwԸn��m���(D�G�)[�%��q�� ��㾘4-�o� �h�/��?Y�E}���IAa
͂���8S��U�@A6��Y����a�|U��������8�~����@:�h���1��Z?���/�I�Gǭ�-��4ˈ����>�`�^M1}�V�o� �B�� �se���&�

��>�|�s����K��]m#�z��K����т�#���5�v'�ڃ(�G�e�OH\	���)���~N���<ӳ&�뇝{�)a�z#-�f ��_�:�@��R�X�K�]�"ɲeߐ���L=�)ߒ|:���݀>�ѯrS�?�˃xs9�����H!���b�#ڂ�����Fq|�DK#��`����Fs�vި�f��%�U"���Dt�Ȝ`�4���[;�`�.�{+�2�Bѻ!G켡��d-.����cHo| ���s����->~���$��,؈[����p��n�1��O�v.��(���.���G�c)�]����������R�Rp�s�US�n(�\YKM��,g��L�Bu���Q8b�g2�̛���ߒ���m:NV3q�x�mm6@�P���W�x��h��U�n��������tW�%7F�h����ۻ��B��M�X7�(�F�}#��:-����Iԋf��<^�jp~�
�H�����s},`R��>��1��ZB��,5C���ag�W��ES�yո-	��K�"�k�.�F�L�K��^9�ƞaP��=f�vߪQ�H�0�\��eE�7��#�sL`�o�4xp����t!��3�kF;��Q�łuFWُC�{��֟X��vL�2�xN�#"0�V�B[��R��Q�[kgX!_d� �;ޖ�+�0�`�'[��p�'�P2���w8vDK$��/<oݏ�mp�$V��x](���o��^N)S��)�g�ӓ1�A�~����Q����w�����öcj� �|��y�QS����2X�W;�
pj��E��t�^U�a$M�ţv)��]��c�XC�V!}G,�r$$u�Z��u�y唔�����#�GI�_�%��/p� B�IW��s*�|�6us璱]&p���L Z��8a��c{����[FVl��U'L���Tr*~c���h��a�F�2�F��g�ih�3�Fa��[`��yB��O��ɺ��%�t3�/���k�X�j�I^-���f�z����X�f��LCz@�b�W������|Gُ7���~G�p囍p*ȿ�U����W���;N_ e���z� �Y�I�K�I��<��W�a*ks]ϡ@��b�����頝�_��7:Ŀݔ�_R[r
��� NPh� �Qz>�M�\N���9:�y�Ъ��eO�M�8'�;��Xq�/D �G�4.}���������d�@'/��֞��#%��h�H'�U��M� <�s��Y�	=;e�׸���d7��tS	�������|��V�(A���,{x �*���!D�,�}�V< �h~ŋh�~�&E�4�I'I�-0� xǘ	T��8�ә-�4�K��j<w"D�*��F����O8Daߕ�v���u�r�fZ؂Y�TC�G
֎+�C�J��y����iux��!N�"ʅ�5���=��W{��K� ���[#��w4�l��Jb`��V����_/���O~kזJ��N}��PǄ?W�G0���^�>ys��7��T��+2gU�x���O��6͠`ǝ�R��.�XĦ2��l�r�V�W�����z(�,���؀U�i?�Չ�3�u�]����<���=����f1� (��Ê��.��dJ����B�L��g�	(W��.��ʧJ/^Y[YF���k@A�$H�D�'Z��]������N��n����J������2�"z�(��p`^�:��i	�{�;e|̻Kf��1�䪀�,`{���w����s�� � ��5�:].�S�#����%qH��k� ���Ƈ��/�T�BE�C�'���^iQ�/D�F��c����Yf���vt�]��2fpw~��	��y&�.�bE�X�@"��ӗ��W",yݝ̈́�L��2vA<�;���.�hB1q�1��)3Y
��{Bw��6�k�.��ir%1/)j�"��+�66%�,3kE:^��~��Mfr����L��<�&���3u	
�U�+���*��݈.#�����4F朳)@C@l�,w�Lj,�:f��gQ�������A����EI�������P�%֦u��f��~B��#b��d�;�'\�M̻.�URF�ą�/v��o#��	FKiJd�4�6@ w����IJ=$��]ٔ������
#��

˯�ǁՋ��N��SU��g�5S�|�"�'��f�~y�"(��r�<f..W��J�G���~;Ј��8CL�C� �Nw�7�c&{� �h�,s ,�;RX�ru@����2r޺�&��uϰr�`�j;�����voO�D[z`֥�v=UA���h;~�!Y.���Uer� ����(��_��WHC=0���U�#}AXYi?�`�;`��q�h�]�-ߠ���I���Mh
����Ma�� �_�3ɖ=L��ȧo�?����h2d3�DI�qb�^A�W���~�p�*8��r;9e�	}��rw�Te��ҸÕA�(Am���k\����G��[oٽ�5V�ߒݣ��;\�4@��~A�4V~`R�E�Nt��L6IogR-�ad`,��F���eA�NU*��G(-m���?�5F�#)j�Z^
="���+o8o��FRŃ�A��|1�e��<�}	ߥCi yݐ3S�[��8?�s8`��kp�2.�.ʴ��� jW_oG�a}q�q��'k+�im��\��9��n��\0M�.O�"}�Nb��7�HW $m��@y ���>2�i�����@�[D������1�<�J
(��aXNl�O�#�l\j�����+���OB��Ň)�{&w&6<}�>;<j:���S:���i+� A ��ƨ��Gt�Ov��li�<+ ������c�����aap�"\��?����O�]���˴�	�*ʖ�<����ݴ��H���h�|Y����}�������ٻ'$p�U-cl9k&>��B��9�s�+ќ����!��̂�aa0�ЩX����iAf��完�gs��mݳ�1˴�V������f�z��n���uS���i�fPk��T��?m�C�����!"H�NW	m�K+�"e��y#�_Y� � j)ǟ�#4�DuN�4�3R+�wu���W��c)6�@��.��$�]�Ƕwՠ��E�����5�"�k���R)�5��]���[A^���V��}?&���@��,X�t�j��\t�IG�G� K���r�%����bԮ�2=L{e��t.�#���%�:&E=���qX����P�絫Zql`1҆�2v½��S��5�4F�jv%{�"⻲Nm|��|��+}V��=pQ�i���g���;��BC=�K�<��8���N���d��fv/]0�)(�)�l�E6��h)(�Ș��s�\�?�%y�%X7����H�{�%����^�92aݲ���b�CV��LƠd��ϒ�M�������x�>��Oa�}�g��Ȕ�3�|xC�%���A\^ѡ�=i=�ϋ����6�!����M��i|ɛBw��u^��cJgid�cQ���b~K���mB�\X����F��<w�1�n%��� ����]Ä��k����Ǩ���"x�@�����9�C�� �[�=̛������f�%"c)��F��D�ܒ�P^�(�	�q�6���n1@����=��ҿ����:�w�$/h��W=.��楻��ULGS҄�}b���O�1�w(\z�2��q��7>����E>~x��T�-��w�a��u�g��j�>��+��Dzq�p��I��Bx��Z;�3���C.j�B�� 
�/Q=ɐ��|�J���8e����M�Г~�K����4?��#��-((��!F���2^d��~����!lMB�9o
L��w8��,������:X�Px-�!#~`��.'�z�.�6d��˩$]�#���n_v�Mu�Ϧ�A��g�0��(� �78��P�0������!�޿ꩂ�WGo�vcUm#�d���Yo�0�Mi���F�H$
�:����\�%:�D��$�&<����zx-� ����v+�{l�jb�g��B��4�M=�`<���_�(�KP�������fZ�	u`7];��)����L'�T�k �7�x��o�%K *𲜪��q^��D�� �u��P�#�5��.�W l����j����\M, '���ʱ�N��<~�4�/cC���}�-����eB�r_�C��x��C������4n�'�w���|_��M̓74o�ϊ%�����������!4���'�7�Z,x���+"d��K�%�|;�����JN��i�[�`����L�YR�)���\���(� ��ꮨ�D��ɲ��d��M�0�[�}���:<o��\ѱ(�忥�	�%S����5���'��� IS׼�:9�>T%1C8���uFf�q�oyE�ߩW"j�1���kN�`}�a��������0�һA��G���gK9��,绪��=Nm�����0��Bo�M�B�9�iI����.��r�
b)�,��s�&8�xO</?��;\����C pfd}c�̧w���*m�� ��#�X�~p�t�?�̕���-u�.-��d����^]ux1c��J8�ZC>>�B�i��cз��H�zp��E�tՕ��e]M��h��l�t�T���۳��v�r[�p��<��WA����
[�W{�b˘wMń�!ݗM7J�mOIf�He��Lf�7���?"d���R��^���ӽ�Ub��>�E�6��rZBv�<��ʠK�p�*��+kzn�"6�r��t	G[��um��f(ULn�+~�m���T�jF<��mb}�İ8�ɝN 4��1�.5ަ�R�k}+{b#�fq_���n�inРա;���i�9M�C�:�~3ju�b�b$�X�_���o�����K�b��0_4���?0���u�TL=�9���bs7H.ڎ���F�*�@�i��s[��r:���E�{ޥ��$$�}�}V��x���oNZBQ��X��٩*�d�[�w;KG��$(CVs�ѹU�0�[ꪮsv�3�6VRԾ&O7��~���D��'q����"ҤJ|�%��#�_H��%���fr�ct�*�:�����<hW�=,�Ly�n��+�S (]�}��Pe{�ښh��E��6��G��6�����^\��W܍�'����Z\�2�yeT���x#&��ϡ�[w���up٩Z͸���
��Y�sP�󑼝�����ڽ�<���T��"z��U^�M~�VQ����!)�9�N��Or����g�|ǝ5"��ʋ\��*tN4l
0y��h+u/�Խ'���CH6��Q�unxˡl��T�N���B�M�\cZu(wG��_����?$��S��ʾ��KKk�/R)��s$�����a�~�E�3J$� MW�'P�ת��C���yK8�E��w��5=��x�]�Bz��>ڏ<Í��TP%�g��y�y��xJ�M܈w		x�r��r��ɀ)�a�YG���P[��e�pһV\]بn�Ŵ�'��b+E9֗�.��@��c��d��'��@!�t��}f2j���tރ�F����N�@Nѥxm�j k��B��S�␡k����t���f�9��x��
�z�ND��[�g$p>��-j*s�������C���&��1k|�7��yMJ�'I�W⚢2���n��×#�,X(����:�et�@%��;��5�[x�m�5C�M��'d:u+(�-f�̤\S�aw��AH�#F�V�ǋ7��|O�la *B_���s�\�	WABN�Z�ڞm1�N�3mm��!/�?_�X�a?�Q'?�!��j�=f�	���!��r~��.N�4m�u;,P��}�ڰ�u����q���(n��i+�8�#������d)�)`��2K����]~ �V�fܕqzOΤ�º�N{���G��ëu'^0���"�FWU��F����9�ā�� �8	���N��3�+�@�uch��%������E�$�98L��d��~w�i��1\T`�,!;'�g�cAϰ���v��^�P��az[��qe��x��qU�a�03�Q:��/ş��K� �4������kc~ͺˡ_q9���]H��{bh�ò7��V��S�T��+�X5������m�d����/M�O�e)���em��S3i�m��fh��.t
�[��^-�݇NU$��I9����D}].���cl�X�N���J+��8�����E��8��w|f;	��ڞ�ߞ�y%dج]9����Ѐ)Mq_)V4�]xU�Z�"��^{K����T!�$$d�QF�ʒ��1��[��\��������]�c87�m.!^�Q
�[�=�Nݞd%ubĨU����S�QP��^k�2L%�+�_��?���mذI���lB��=�<=�������!#c��e�#L����v�L�gO]�={��H���H	�H��L�fB�I�Ј�B��m����Efי �b����']�]�01��a~&���Y'���9��U�Zh���*v7;�j&<L,�ؿV��NW$>2�Ϊ\��q*5�kJ��G����4�D�ɲ����KY�k�jg_�LQ�}�,݅�l{F��X�6�!{X�9Eb���A���A�K"���0�E�9���B��F�a�|��#kD�T� �C�����[2�jE������,s�l�Od�=��#�\�Um���k�{�W~z+
�W)S�䑙J��R�V�`�I>Yؙ#���t�CM����A�*F��S�qy9�<V��������.��b� ���}��ɤ|����m�cH�{@.D�٠���W�B���@�q�����8�mny�1�hSE��@{�%��WƝ>���׏j�Νi �#��3�����
�5����޻�:����>rQ��		�E����6q#�є�E��o:S?
0����@n�_�S��B[�+ĩl�|�p�Z�i�*Xdc������w�d�k�寇xH!`�[H��/>_o���V��$�2����4 ��cg��U���UvqttȻ�Nx�k��!��@1����4������Wh�������l!�^<����$��SEe��]�(@3�'������5o����0�w8�IҶ]��V6���n!5�����G�Y3�nr?3��8�LQXKw����+�D�3}2��4.M(��fD&ˀ�N�l��K�	-f�6���M�x���(2#߻�������1Y3�ш����Z�R#v���V�*�q��w���QV���PiX�l�^��^���d��j\(�_�JÄ��IQ��H%/�S���;	Y��s���m{���D�'����8�"����wp8,S�S�w�z�,�_=#W޷PI�*;zo�朒�G����f	)��������#lh�d8^b�ɽ�5t���b(���)w�:u2�d�7�8�Q�P�A�,5K���e��ϭ��I��ہ��q�zv2z�'|�,k��b�f2���6�b�^�bK�É5�q��Wm.2i!���� �������L2���W6�i���~�p�we�(��2�.�3 QSk��$�/��kQ�2��@�)��WY=x�U]v�=�DF{	iL�5�EH_�ڂJ5.�D{�d�ܧ��57.�\��)��e�|pSn��ў�/U�1��DsZl����7�Fz-����gV����Az��F��\:��@ߐ�8�,K\����	�(a^�� �d�!ɋ��cd�Ҙ6��N�|=�\5!d
+��ʳf{<��lf��/��Y<�Ag:�r�嚊h%|�:Y�ld#N���K��t,��F���s��l���p<DQ�ke�<�y^��%�+��%�X ȕ�M�+2Ӌ�O:!�#y������#U��w��w�*�c.#Ɋbs$�� �Lm�B���&^p/(뀗��/�M2�²4���	.�ո-hU_i�u����P��K<�2#����X�x{���HO������s\�%2�$�����17�a\`f����2��T����$@MP%(����gw7R6��װ�gZn�v��/��\��;J����i ����q3��6�'���Y˶�p�+1�\զ�a'>��m�ц1.oo9�� ��E�F��I�J���"l��j����[_ż�7+;4�V4&q=�{���e�+��xt�E�p���V�������4�;�R��S�_c%�X����̝�Y:6�C�D���VmmU"Ȃ���T���5-�2�����z��f43va.Ztei�{�섁.�'4O��'�r^��0��Q6S��*�q��t~oAU=��&�R�48�+�=)�+cfgR ��I}7�r���@���iKq����
�;�����=�Ѥ�K~H���5Y��u�A&�g�b)��B=�ٽt<A�^Jx�+��W0+
C=���z���w���U��� <֠5gpm��K~aqi�Σ�S��b_V�'fgJcM�B��)G��b}u��8��<^��	Z���Im�i���7Q^�׊�U��'eg���p%��(�ۻ�e���� S���M���g���uP7�(j݂1C���#&�^-UJMa-���a_�J���&�a�j���$��˸���k�vxꏦS�9����&v�F�΁�%�/� i��O M��_�/���%�W9#p����u_Ȇ�����7�v�)�m�&�K�+ ���>wKF��YN�ҹ��$UKshe�����|4�A�|���qF��aO%���Q����*���sըB5P�����١kt���JxV�'h�-/�ˢΌ8-���Y8�*z�#���˹�}W�a��#�6Zw��$>�D,R0�h��A�-9÷�\��^U��OC@�[v�<�������Pe�|YU���:��w~��Vҷ�=�=��XúG�!��ސ����>�([�~�@�حۦ'�.xs�&
1 q�$�'P�g��HTT��B�[;|W���̲��A��v��ݽ7���"�`۲�,�&߽���hN�έ�޺H�fƓ�uj�5~��}���ܼK��G,	d;����W��nH�I�t/����+ a�^�
'�ϙ/��.��񷨦8�p�F�̻��l�fA/�`Vݵ:�J�';/���d.���/c�Y��4�W5�:����0�o8_�"E�@|su�o9Զ`6�[��R���ہ�	���c�jK����$�D-�2`���;�S��T0�A�"-�?Xy0���z>o���U-�ͯ��2��+t"�(ٗS���?�X�;�)�4��g�!�a��h糉l�O|�����#��YQt�7rtl�'�RB|G����^˱���]-7f�EkG��� �\��N�ﱖnC=����k�ڵY��Za �v�a�G�.P*^<^#���i�̚��P�(�e�n�`)��O�D�,���p�����߾��V��<����Ht%��7�����{zC�����'ː��L@R�pcZ�H[�M���ܢ*�)�����ȅ��[����rf�#\D���P[v�9M`yA�ޕ~�]��Hb}��;D���#�����J��rce�A�#���P���4���Z�7V�䅯/4(�!�W�"�W$7a�P6=��0�)��x���?+�A�(����O���a}��}�9	Q����p��C�� ���,YW۪�Ц"1�8�]՝�<��n��>��S���s�3ϊ��z_T���t\_�QJ�7Mɡc�	!ٖ5��ٯJ��3+Z�h��׵D7>@Gͤ�j��
��2 ^�����H�Y�k�q��Ɇ����~?����[#յ�N:,�A���V�UN��YTTg)�14�H�3.��E*�e�Э!��]R�ڎ_fKcv�!�Xb2�O�H��>���+���a[R��BW���+�����D�~�tU_��6��/�1F�N_m1/A�4o��J�F��,w�c�bR1��Ց��cC��Wm�[E˂�Ro�Aw�b`~�r�B�U�����4*d���&�?\�2L�4m�]�����
�0�K�'�����[��x?�x�\88Y�\�<, G������D��(�')���o9k�as�H@�LI�®� ���m^�s������|�2m^��^R�P{Ui�����P�6���ْ{~� �Z���d;�r?#*�dKX�A�\��`5�	mx���1�G�4�ǰg�-����5�/��]��coWS��&ćC3�?��1*��F������^��e4E�,�T�Y�5?�|����bv�Z�zv�j�l8lt���$���mNd��݆��p�"�ha�>��^������۰q_�r�\<RC����`��frP�.���Y�rƳ�f2�����y��_�?9n�뛞��@�Ր�-��B�g���{�<�Z	7Y�*�_���*���R_%�
Cl�1�>�3O�s�$�|�N�fS��얺�U�� <"�^p�B����+Ņ����#�~�f)]�n�>�p;�G^^C��B��#�a����T\�XP���~v�X$��c�����|�u��{ͿXY4�)�'�G��5vt�����>�l<nr�û�j�ȧ|�0��ժ̀%��Q<_pKS�wg�M�;�<�<g�ɜ��(�f���P XY��t��ġ��U"�hԼ�|&�d��H�+�V��wF�@寂uEJ���ؘ|��b#=�'��0����	�$�X5��a�>�[mu���)џ:���	_Y1����P�ãmie=����?�����r����"ӽ.�I��Ă}�r<&���}?O��.���ަGI��Z��C,� �����Ić��O^���춍H�D�wbΚ�<]���\@��,�y}~ކ��}lI��u]�2�޴��)(�O���s%8���O�kv��rbPp~s��`�0\�����[���}�Q�nL�Y�2��RQ�i���$ފ�Mq�� #���.���6�2�4΀���V��uI	�B[�o[_nU�i����5�X*�0þ7����B�R�>kdZ�c�]k���t�n:q��%���N��r1{\�E�EFl���5���i#�܍��c�!�)���2m��!Ѕ��sЄ���,�[&KC	�qWx[Ua|����6���<�^���g{,RB{V�cN(TK�P��s&v�������:ߜ��PC��������ս^�I%�A�n�3E�n��7D��4�{]�z��,��P�Y�m|ĵ�&�m�z���#�73����N;��iu�D�JD�+�E6uͅp�$:�����PK��Fc���)Zڞ|?7@*�|�w�����L߄Old�̶�\��?�{��ՆA�hj�����_���(�����Ԛ`5Ou$揼�+�K��"c������L��W1LK�~�I�͂�nG��N�X]��N�=�F����U�z�zL�FP�[o�SX�Z��/���|�;г��h�0��Ldg��}��'�"�wC��q}��tDy�U/2W�>�✒b�s$֟4^v�{е���uS7�4�j+/�@�[1�	��}CG�7�I�I���"�qR��������EӐ^�Ъ;%�G-��NNbÐ��,�ls��@�I�A���������A���'�-����ٌ�
�ᤌh�'E��R�K�r8Yɫ(��2;�0%�Xk�w-�>70$�x�*���۴G���5>��R�f�{��K������?��i-��i
�g�n"tlЊ,���G!��Í�D�ydm�h:���h�}�z+�����mj�f�b��j
�7����!��,T,c~�`����o��H��QK��D7tu����GC\��Td�?K}ΉR�/�
蚝�c������9�5T�'YR�Nzyi>3��8cT�³V����eam.`08Օ,�w3�mq�|:"\�_QCR��+�8�ݠi�U�
�W�NG��(������v�Ů�:AK_�~�%���K���@������4���~�a�_M����̚X.�I/���y����`D�JLê���$�`8c����,ޘ��"��AS��]O�������m;����kh���z=su��s��s�o/c�7R,7�c.!Q��b1���(�!�Y���H��p�s�z9�(I�\��-
??Ok&��)�f�HZA-�O��a�H���ӆ)J�9F��;�)�cf�oU]�g`4#(��#�T��yS��ߑ�)Z�>U8�Y�p��u��}]�{�gb�^,l�O�,/q�4�(v��兕NL������jf��KWlz�i�7Kn��T���`,��v�w�����?{����F�$JT��!}>U5���bY%a�p�U���|��I��?-�}V�<�Z*t���k��K��+�$��!D�T����3}�ō\�KJ�*��t����J�S6���34(��(��Z+�s��Ll�8v�-D\�3�-��y�xc �j�*vc����͚�q�֎�1��4��ŋ?�[)�>	��׍⥨�CVՄ��
�a����k�UR]��8-%e�R}��y�)����Q1��r�}隣��$I#�7Qhڔs_ ���؀ӲD)_�H����2p���@�>TK4Y��Ɨ��&4�%䊑B�
��2��ko��a,Uܡ���L��HL���~9.�в�h2�g"=��H��1�B5�7\�K/3C޲� $%w�mm��+&�#���kH@��m�3\��!O���α[d��4rZC�a��(z��e����:|+�;�C*���7�;Ґb`�Yϫ�Ɛ�0��F���C� �ߝ{xu	��H�*���E?��%�r��������@V��L�)���nL��,r��5G��oL��B�߹���W��=�O������,5�g�g|UёJ}�C����<���]j�|tmz�W)�!��X����b��q��`��K_�/T����9�'��?��������?6Ԏ���h%F_#��J{��@�m�H�b�Y0�ciV[��c����s�:.0�eu������j9ۣf{Ȩwn�3O�7�*��n�|Ѵ�J�~�0J��)i�	~��FU�v"��[�e3��&v���������m�--Xx=�>�J���wh����a��<h���]��Lϝ�vT!aF3��A�]���Ta*xLU�ԚyU�5���G�̘��F3�W�(���l3�X�m��Dڶ�{�~�S��2�#8��]�ф,p6q̺�JE��F̧9��n4��PIf����-���&q��X:u���`K(���-���2�|1���%Z�]����tPD�u���N���Q�݉�����N�W8>+�+uv7�V������yA���'��	O=�%�2��!��lS�㧌�	hS���0�64'��j��;��f%24<��~ ��"?�F&�2�m����ƈ��@ɰ~���|'�PsX��P��R���Eܑq�d0�0=?	r@��"��Z��it�����z�M~1�q�;+�8�G�D�tڒ�k�3��ᶥ_������L��(��9y9C�}`	�} �@�����?�G���(
ƷA��=�Vj��pGr��_��מ�+F�FE{k�L���qJpBX�iE�x���ۘM�Z��2ݔ�	ܵ���[�瀁�A�ϓ6t`h��7g/uX��E��#P_�4����TF;!�(W�����	p��e�_����=��{��]���{^�_'uO�#�p𣈿���zU�oZ�˦D��nU�T�\�~Ҹ�s�)����l������Rٹ"���yi'�y_�0�ݲ�0�^c���~�K��)�N=�
�t)�n�F�ੂS�D�K73.�XA�8_�^�g��ZQ��_��r�����L� �{yk���q�q�<D�9S7rlmT˔��yߚZ���� b�[������\��������J"��}�P`�~�	tY��O;}-�\VB ��C����e�e�l&��ksbN�������lj��Jă�nr��>��6��=���ƥ��i��D'iD��"��D�(��_�ɬ��Rr �Bũ��\�
ms�����cXڄ>/C{�R@�v�;ek�*���"�/�ң(��gP��ٙ����7*��X�$����__��ݮ8ޞ�����h'c�'�T�)��rd�a@F��0�[��z&fM����
Yt_�������t3X�壮�Ѓ8_ڴO��<?���Ι��u�Qy���	���z����H��qJ `D�����F�6½�܍ϕj,΋��ﲕ�;�n/l�Q�0���O��}���,|��aD�4��Q�R%z/�0��U�nL�E��v(ڒ ����J�o+F�ﱥ̛��<�Zx�v	���	�LYA_��Tˬ
�/�űڹ'���
�Vp�O�Ő�y"=>���'�tR�W\����@^ljr�e ��`�����s�S�����I{z�wUy��|&s���1�j���PE_lK�)@��F�t�Q���������J��(X˒�@��9�̓�aK�n%5zl^�i�۴�+;����PiԐ<�=���^}M��J���,����9��_ᝊ��:K��j�>_������TS���]�um f?@��3��. j�~�3���4B5�;m��"I���#R.W�oO���$�7�����2����`d���0u��n���PLv4��_*8`Bf��1�/#��i��2v/�%��rNǛt�S�cGE)6r�<3i�2p��p��D���_��1�V�xG�K�y���[_��bx^�a����9h��B��V�;���ALR��.��U��u6��51KBR>�j�Q��o��|T��"��3��!Ě�c����g����6k�+%�_y��j�e PNHK�/�$9�TE�}He�KMsqڝ1�w��R�wY�gb�#q��0u��f�'=�\|c�r>�ʷ�ح��M�E]���n\)�x�:��5*CFw�q���_�'*�.��>�6�A��F���n��D������y4(���m��M*�Sn/EYW?�d� �RaJL�r��oi�\&�	4\L�����G�J�8�U
@}�3BE�[�N������v:%lӥ��/|�hG�b8���9��P��a�Ŝ��{�·�A�i$&�'#� l�>��*����gn��� ��nGް�~�/5�=��C*"���n[�w��М�V3�)��~����C[������BP o�R~��ABL��뚄����^��z���M3N
��n�е~�Фg#������% ���X��W�+�2gކ���X�-t�W�+���}|ν;��]�>`�ǆ�hZ[����\��P�L-� ��4�t ��K>�Pp��;^����U�,�N}��$I����s�a���Fш�?`h`���c?����0m��8�j���a8&^��G�J7r�f<�a���\�IbxI�qD�$���>0�ٛ��gZ��pǭ��=��.]�����.Z��<O$�	�T �EtX�ۜ�h0�3��� 81.̒'��G����%>��F�"!�Wv(�����ñ�I�ʳT�!��i����Pg}�Z8�� �H�B�Y��_d��	P�ߕꢚ-F�-�<ɦ�:�Y;P�DoF��B1�C_�B��aB���:>������u�AQ�i�x5.���n��)(1�6�Ĉ�@6��ri6S�?ޣ~E
�����ʘ.��:	�M�dC��>���"x�4�LG�����P�#��[�O<e�s�"�ڮGX���o��qx|+�5�o���ݺsR�L��(h|i�j����T��ű���F\���!��Q_��n�˂�n�r�gL+�T��b��n%�����9ix�M��kKf^� �Nat��H��??�pTRD�XW��j�0�i�.%��մ�:R!�I��U��c�������5��ca�gf�$�	��-���+M�3���K0��y�z��������ͩ*'��46��P��� 0��@�s�H!Z8$��K�M�獬�P�Y��}!;neo��VZe2ZG�Ǭ���-����R��I�	��'�����ε����≽ZH���"��L����8� [��;��u�h��~Ȍ4a��`h��h��V���r�x�'eРW
)��&���,���{�X_˖u0� .��J��L��`�ϲG�y���J`����c�:�K���̛	t���v3���~;����ߏH!�Hѷ��#FD
w�b��lKY,�9��	��t�l{|Ʒ)BL��w��X�ny�F��£Hq��i(�A����Z�3���f��=�e��͐��7��=f��]�0."A�/lX�O�L?ۧ�Ha'/\������;�/�+�@��'�CZ�~CˍK�W*�ϗ�#@>�k�WD*�,r�� k�!���,gt��ˠ���x@^��t}�gkE�����^8�d���"��S��^Ћ����
���0��QW5����*��V`:�CZXu8.�
�1V햄�_O>�u��J�_Y�:�W�1՞��4Q�HD�.j�O�J�RZl2u�N��L,��ʞ��fh!��s��iZ�)ۛ�ߗOGW�<�����ϝ|�P��g�`��bn�p��?y Br�,9������YWd�Y��9꫻vԛ�Le`�����Z(P��w�ٍ�᠌�g[�1��xP�9j��JzN�^9�~g��k�Ȯ� =s��j��8�:�9��A�T���L��xߏ�Є�[	P�_�X೫{Y��^��n.���t�.~�$�</-�=�N�]>��jkZ�
?��p�a�`�����W#E�W���#u�W�!� n�bv	X����A��А��bI�@�e��XpwC�j�h/�U%j|HDj��sn��9BJ݁�������<�Ź`�_a���������&��l�R*���u,�t�T;خSph$N �mˁ�J�ʺj����r���=W|ޟM5��P�c���\Ym�)!�n�E��U�w529���Ϡ�y1~�D��Ⴖ�me�rk'�����������Y�>B��%Ay#�=���~�ψ<�G	�r��}�R/��p��lz,C���OY���A�y�Au����h��cukB��0���ݼ�����3��m����U�ܝEptp����ez/I�3�CUE���bǗx+Yi��}�����ֻ�W6Tke%������)�"͚/��~�w���hGu���$��0�euw~L[G��˾n��p��-��g�8�:Y`-�O�������x������J�i��}���2��o�h� �Ϧ��pq]��@}�'�&�3�a�bR0z�M�aűh��@U���{Cn�:�]��y�a~Z[���h5Y�/	��otG4�Xr�^;6a;̘�	���`w�m)^�G�O��-��B�%�.=�q�o�NV�ԇ|��R���E�=�э���L��bZ��AY@�
\�+�$RT��Pp�P��3H���@�|ʺw�@��>�Iq�%��Y����)�lb`�$��<Mt�~�j�U�j�B+X&���%�*��=B�\y�է,Ki@�?��ҥ��$���-�ҫ�n��j�,���7ۺĖ�H�,� � %�GucTPGt*��E�j*�z{ޖ4�uAfY�jU�?}d	c�� �=,͊�yu?�*%��Zc�r2q�\E��g_D @�/J�m�G��Ň*k>�����%Y5?���
K<��XL4�k�`��?�q�`G���� I�>V�]� ٸb�&3t�)M��(,3���D�Kj��$�cZ���W*P�q��8�R�()b�.�"ŸA
�� �J��@�H3wdyq�n�T���F#H�n$� 5��V�<-g��b14�4h�m�{[�cl�,��G+�'��n�D�8S`�����oIxn!�i����������������M?��؍��0��g�ں&�N���e�ܛjNЎR����N0������#@j#���EU`�78�r'���y|��GO�)0&o�v^x�ؖ0�Xw���V�̻"���˺�Y ��y#M�Ey$��
�ل�X�@Uy������=��04�d��D��1���ɤ�.l/���h��X�SCF��5/"p�g���6�c����IDe�R���ݭ��$��Uj���S��fD�f��^R����:�bѓ�of���!׺`3g96�7.�tw%�/*{��|��m�X�ǳl�6V/4�ޯY� 4&���S9���=a���4�15-7�$˗���%
�l�D���-X��A��mS�W���)L�����М������5jR�J�r�A%��Cm��-����٢?
�7!�:�w��Y
�z��J
T�w(_yEk�?�E ͨ׿M�CE��������U��$a�-���/����%��h�c�R�� N#d�`^>�ǿ�1�@~#��ZBk�N���0:�:�۟�7�?p�O9N�p���KwD�����^ ��"�9�V�'ɳ���#���*�~I M��Gz7��mK��5i���)$���/ͭ$R�A� ��6[���Fp��S�r9�}+�S,�uPBb�L��09˩5��q��=s��ë�5\-z�1�uU�(lؠ�8�ɘ4����bvC�s��zc�$�s�(�lzZܝ�&�*+D�'֎���%��*���/���lel�Z�4�J �����q��6�*���|ůvK<4X���WpOD��7W���*�C~��y��,<8m�aZ�Ĥ�݉?zX�'��5��P3a�U�iO_u5\�&�,�!���\�F�y����G�4����k�xq�����l�͉�R�{�a7ÄόKB�A]�ԍU��X����^�S$�(��Ls@`��hq��[�/;L:����5y���D/�2>����[�D//�+�@���))�����8S��X�ģ���e�"\Ҝ�B�s�~���x��ϛ�ĕn��G�V PC�L�2�+~��:�g3K����~Z��V�(��D�%��/؃�f����rsɫ�+&��z��Z�O�qxZP��؄���{���KL�̸%�@ݣ~%J�A&|��°�f%��尋4��Bõi���d�z���9pA�LĈ��J՘�.h�(j;�Mϩ%��Aw�Kf�ί,'�փQ"_P~?��ޘ�.1j��C��W�S/���{?�p��"�^�znG��^7���ʆ��c���ƍu`�!�}=|�;y��M�f��NلFJ�a>�V뙲��˷�>]�V�"L��넚Ű�Ȓ�{\�v@�Q���<==���oA-A�тj*4�k4N�K���m����K!* �הǯ�Q�Э�r��9�)�l��L���
^B��T7�9a��3"Kx�����p0�=�~�[�"2��1P�W�p;�`�f9�	yHq���]�a�@y�4�����e��f�D�}4�kz��� ���;˂���ݕ9�e]u�Y%��v�(��r�h�5 o�A�0lb�y�̱d�q�7F7u�L[�v��e%V���
�l���Da+��݈-��>���E�=�Du#���!*d��R��E�����0�Yy�l�װJ
B�hN��[Y�X}Z;W�P�C�j&]&��w��zvd�����[\�21@8��{zÅ���C��i� �ha2��tm�1��y�"uZˀ�ZZ��m"m��ٮ�5lC�.�HC��{Y���aP2'w��БI�$�//mX��2�Fߞt�#ec�4}'�X�Ah���� ��8��y�>>\�OǑǳ�z��Y�u}fY��6�K���(��ɪ~��t��$����N�J�*�ˠ�k�|v�	���#$�C^Ȗ�ݻ<�B��:�C#[2��
�R�'���a�7�'[�\yy�'}�->Yy�Xx+h��6B\�i=g7_�]�4}G,HiRH�0����vx�q�2b�G������ӧ�X�eq�M-�}��&�����
�E���>J��¹��1��y���^��\���v�D�#�$/viI���X�,���2Y�l�a�s8Ѹ4��D�1�HI�x ����u���*ś+:���W�Q�C�����~+� &��R��fmd[op��ƻ��Ó�U��U/ ���[�n;�Ţ���p_�q9
ݎ c�E��u��$���4L��h�H��� ��Eҍ�"38��7$�*dڮ�"pva�8�!pC�$̥s�a۱A�����- �Ⱦ��#��c����'ޓ����/�_�<-�)<�nW!pݛ��	���Smݩa^��8qߛ�弉Fd��������r�U�gpL@b�Δ
�k�F�R}Wصr;�M���{��v�(πq����qbW�ooz������[	��e���,Ͼ��B��r1���Ľ]"[�'5Ɯ-����z�/�B�^J( _#�N�~�)z� j��s�#�W�T,�H�H���|}5N~t�.�^��%r����up�'�8�5��U�Ly�H��]�U~T�YcDo�M{en��;�؅	9�mӂ�}q�<�D(q6/�)��7~v�f��z �2�Ĭ�~+\��2L��r��ǋj�;I*��ڋZ�'���W�P4�B7p1CV5�B�����b S�Q�z4Ƭn��W�06G��t��	���Ȇ�XҰ���<��jժK��ʩ+���C�L��>�$f��8w����L�0��X�y���!ǅ��i��\�w��/�asA'�bRt��5�h;)�����Y�!x,�����y�i���q���Ί��}>qi8�gLq�=Go��uBRxkN�m�Q#�!S�e�`�ĴJ𥥍��e3SV�
T��@.���;�ߍnF�M��B�9�IAE�[�@)n�o�Y���%<7&�I��d��	j�&̀r�$4��dr�N����^��} ��!�M���Yt�P�z��m�Σ�r�􇊉L$�V���1�p��!K�ֆ��
���R/�ǁ#�X��0{��̀��`n{�sn�F�3)��y$ZQu�6�1A��"@ge�l���?f�����G���覭��O4P#˙q���7��}��?��?b��7hJ^
�Q]�@��&z)��J`��O�}�\'�#p�B�[�8���Z�Ƶ߀v������#$,��yA��H>�O��x���y��$�mm]q���tG'�@=�"�K}�~F����Ȥ0�G���������J�6Y0���T���;~_L�;���쫀�թ�	��c��G����Q@���I!,���̥���;Y���5�)lwۿTv-�صҕ *�CR��p�>)p��H�������ZE���T	�3S&�xj@�kT��~��H�m8�z�ްj>^��mv��-���a�K��� ���^/7'8�7��s����&a�*�{����3��^���l�ٗ�mq
���m���29�mݧNd+AK]�%)�@������@&}�G���V��Hx�Е�a��~�~PV�/�XY0���G�w��LR-�]7��CbB;�g$���܎㏚?��ONp4 ��p
(ӆh����'"�Z�|B�)	]Yx�<b9�� ��.���<�m�R�S�;���=D�3�ǿh�:���	�-�!��!���)�-f*�#�lS)p˗�wU��/�o&F� ���`��]5�.�ə�>:O�!U]�J�����(��)\p���ʏ4�g�'���.�Ƣ`�Y k=����}�^��9X��t2��-8@@�5�����
Ē�G��D\<҅ĕJ�a�fSSzp�5�WAY�,��t�V^��6�w�tz6��OY	s^�U��L5���S�IT���ݛ=�yv�
w��bp��d<24���,c~5�tzĶN�w�x�rs�Q;X�g�X�	�y��q����϶LK9V =����:`�P�y�9~��-�;����S�(}��H8�u�]�a���g�^�+Ӝ�5�"{��&����m4�	��nq��٤0R�6�c���H��Z�����	�a����P�(B(fT��
<շĿ���ݒ�E�G�nJC�����H�o(%F���	��V]z�뇇G�E�����T���k�h��
���v��>��Mv�#ۂc��|�ɉu����o=�ض.��q���_��9+yK� �*#d_Q7�dѝ�88���sQ����i����V&29҉.�#�����ѹ�TO{��p,f��/V�յbK}h!{p��T���τ���\L2Pu���dq�K�g}�Ɣ�(��lzF,���PD�|��2>0�`�ox�(���������V0��{�G��I�ٽ���ZǊ	�@~��u��wnA�\F���#��qB���/���@�]Ļ �O���l�B��І�H���3�ف��?�B�;��:��5�-#i>�/�ƀ�hf�����Io��VIԈ��]��
|�G�D��"sX��Q��5w�Ne��X�UQ�0��GA�(rJf0S'����f�[9�l�>����r
{�{Q%Ax��g����_��aX]��5�j��+$[q5�/$�*"ENQ���M�����\�2V��:�h�̙\S]��'2zЕ(��l���wy����dj��ۣ�@w����[��yV�	�zdk�R	�l�3��c�����Y�wn�Ǧު����1��� �b�(���н�+hS�����w��[-��iY��U0���.���(U6{
cƵ�x1@��Ȳ�y��Th^<ˡT	���{'�<�|���ޭ��_P)����_h�t�tm$���}��7Pp!k)7
����U�3�4�y��	�ѝ>�ٔ�P!OPe�ȯ2�t���D��n'f�:�h�ΆU��7E�s���!T�'��n��,el3&��+f߰��F
yCB;$��ɓ��c���
��v�|ZR-�x��0ݨr�{Uh�9dp���|Q~�n���8�ҿ��+�#�f��_�-�Ӳwɯ��䱏��zh��O-V�'�-5P��;��W� ���b��������sUo�iw����Ko�+	p�w7b� ��?�@�Y�����i?3ߕ��
�6A���$����F�%�G��,����3�bY&�,�;J.3����w?X���49@&���#���Kܣ*಑���1�lS�H�\KCj�\	D�8ck�Hc.&� ��;+���##څ��S��+�ф~� |ΛNM��^RX�O4��33���0g2=��;]�#7���`�;�tys|�0�D��%1�wa)0�0P�Xgo��6�����M�y���h�;�����j�qq�J�g�(��$�e�5�Ⱦ�L�X=�"C� UR�l�
2���jX���
�w��r'����Ƣ�� t�0���yf,b�h;�����q�s�^�d����⬘�S�g�J�\'�9Ys�����,P����5q#'�/i�4���$�d h�R�ZJm]
i?�M�%u����-��a��?,�CLv��g�(b�ɦ��M�Ѕ1�Y=���|�$r�;"�tS�XN�p}A��P�X��L�IO��� jq��,GyP�~,�"�W������p���	���^�m�=�K�H�Z��-n;\��(��l�u���y��<�q�q�;�{H��̍lٰD���"��M7-�$P��k�ìd� T����[I+��txu�p�dA��\V	�y��k���+�秮;X��u�7������-W?J�P�x�|D�H|�<�@��#�T}�ԑ͢�aQ�y��׊bܬ7�>.\^�t���[/���F�4��II�^w�JRf�uܐJ�H�O1U%FF�ї&���3�x!�hJ��s�]ܰ�s�!�~���n[��<$������ƅ4�������R(�sԼ�4�h��w+�����慑�	\$�����i��FUoV1[f���v�ĳQ=40����ܻ�"S�áw[[�(��3+��	,�04Q�x��Op�[�O�Y����ë��'�盒!ku㞜�3�8�* �
����&��co�&�SX��`tK
B*�p�Y�V�����@�vK�����"��d�1ʷx	FB���;t
�\�\�!^\��E�ϒ
[K�G9�})�N{����'"0G��FE� V���� I��?��Hl�c"�˂�C^�i�~�.�l!�+�)��c�+��;�e�����a1D��w<����4�GkZp���Z�ޖ�N�C�q��Τ���nU���jUr��� �����X��+-�F+��ǥq�e���Ȫe2_��t6�|��㏦�\Q6[�RQ�Yg2���V�٘od2&���.A�Y=�}��N۴c<<�bC��ֻcP:59�3��3?H�׷��C)�m��e<�^ I�0R�i�xF�0����lL������V�׫�N�N�択����P��2���6���}�?�~�����7��h�Q���7� ��!��oE�O~M�/�광陦M�?�����%H-q�x��(# �F��Gʼ����ϮWWs�z��Vap�0������G뱋��5�)?�o#�q��!���s%�l�}i�S�	�eJd�?�9Ee���\_|a�Z'C�
�6�G �w�a��X5��1Rg*�X����".鼫��B�̒���=o���,�y��~��J�^�}��<An�O�Ui�4�0�{z�4�]4�N�i�^2ƈJ�;E�h�IO�#Gu�����;�ž!��Y�,�Ti� s_�m�����n�qv1EE��E�5^e���st�%ޔ=m�z2���)i�/��M�,��g�=k�һ���J��䮪��zz*��r(�$%K>(*����8�m��T���5�i�]?�CC��@Ϭw�-��<�Hl�}O��VI�t�]��.}��\�7����&�]�H�D�͙�o`+�e���Dݚ1�(�B�u�tW�;y�]ʢ��M��Mt�Am;b��Βοf����%���/Ň�l�˥Vp�Dl��J�+j�4��s�@_��}17J4-D"I.拪d���G��l�.d,j�e��,�.~���I٠C�ݏ�kr�\'Q�T��.(]Ɋ���@o�d��d�~L[is�cy�ð�n��ݹ9ǆ%<��x4U/���J�@��e�C��`�X��s@���W�������_Y���`߯?����\�
c<�/��W�N{7��W�XŬ�jN�ps�7��r��#�G�J!V`ڬ��jr)/'�0tѬX*á#��g� c�l,
EK���y��UaVX]N2���og�=#�pA��hܤ/���Y^[s^�����m�T*�=Q7�p���7�<��h��1�x��-?u�a��h���E���HM+	�g�j���P��j�X�-�ϛ[�ksKJ�-�z%�&��@j�e�
�_���/.I�T~6�P��%�l�+[C{��9�7�{VL"�Q2���H������ؼ�j�J����wZ~����4?I-2��r���4G�"���DiG�q���y��:��u�4ǣ��\H]��I粦n���c��U��9p������=�¦k:h��y\��0���)��]mIeڒl�~�#O���#�.X#�(�fA�x�� jl���a���H�s�\y���n�G,�n�$a�I��HvY��J���
�GFw�Km'�`)t4�
�a�puF��yN?�:�b-H�'v�$f�� �����6U�O��	S���}�g�n��+�	)��o%�=���-�@Bw�XJRnBj�R��s�����1�R��t��r��C��H*2����(V
:2���}��#��^��
��vS·F��8z����z��6炉[B��x1��qm��\�H�-��E��Daƈ{�q�j�L����B�qt֕�F��M��H��7��)���-���Y�!M���V<ɽ��m�tT��77�+���|.�|�T<�V�^���hYE�q��.�C��gD��E?��Z!�]'&e^��e�R����|e�Jߎ�o8�tRVe���ݰՅU"9�`g������xn[��� ��4����-z��ŏ����v�Rhr�+n��g���P*�A�� ��"�׎"*M��I�O��:Dጳ�-,�xv��Δ��>����!;�NKT��~&|b��`��^S�9��V���Hۇ���7���O��NG9��y�ms�C��Qr��;�u���k��a�������,eN�Hmm���{���ƺ��(_��V�0�Q���k4q�m�W�׌�$��*V�/\�$iO�J����Fx��쑲Ӧ��N(�Ճ��d����V�8�4�V��x�\0j���Zѓb�;\]p�����	Hy|�l��C�ƈw(� b���\���~�)�b�}^�:�4���:��_�^·\ \lyV�}� ���.��ކ���B񸈄J��?TJ�V��ٲ���<J�!C�v��I�3��d�/ɟ��0���6T�����)��]�@s��"�X@������I��(aڐ{�4˜(ܠ�u9 �2`fx��[�,��q� 諺[�@����[�>�gu?�&�5�O�߫��Uo4D%��Nl��C�n}�-�	��ߏ����Rku�}��r�z<�['���1)�g�+̈́��>�57���a�b�З�-��B��2AM�^$�8)�z�F-z�0�ޠ�&ɨ�����|�Y���[A��	�5��U�tpF^۩������"�섁�K����
'�s��1Y{��#��M��]��F��Aq�1<����iP�*�����J+���b���D�������FQD���I���}�w��V���S�7̝8���J�lf�IRXN��2�L�Z`��Q��B��z���`��"3ڷ��aK�
�s�H[���%eْLy�D�߭Nǹ#=z^uN3���r����rfR0O��hL.@���~�S>.��͔��ݥ��[?�(D��0T��� �Rݾ~�0@q�Od�]�(�jh����3`���k����|j�`?����&�=��=��D��L�Y�F!+~��`�LɃ��K�yc>p��:���w�aP�@���Y}���nƯB��U�}��>ߎp �,`@CM2b_���<Q�՚�I���t�R`��C��)���2�
m��=�|�<^#]����o'r�-=Hf�d�ɐQK5~=� �Ku�᫰���:ӽ|:� �OLJ�N'��̸>W�wINUQ���ײ�.�:_��h,D+��BMk=�*|��K��B������v1H$JÞ��+��fe�9��3mڻ�&���CCZL�u�QR^&G��"9vN{J�K�Wj�V}���@B��ڡC�|k�Edh��$�kQt�L������u�:��u;��=8�&v��D�lк��v�:��wK���(����RIK3�ŵ��LǸ��3dΥS>��&�Fᕦ"�V?	؟,VU��z��^L˾i���� ��0b��	6��hqP�l)q�g˦['] So̙@��@6m��f�lSmc����5aa֎�*JM�q�������+w��ۼ����N4��0�eU%)wV��n�]sK���J,��.�b>�t��Sn����fLaS�Q��&~����e�.��~�8��	L��Y���Af� ��n�ƴ�9O��c݈فCR׊	�m�p�a*Ė$��{����@�i��@�O}4U���K��8M�2|�l��(�c40U�\���:�j�(	J |L�b�r�'e�������)w�'���x?�r��O&J��3^6���(LY*����Y���L<8��4��,�Ꮻ�����N�׎u���X���R�P17�pA(��D���q��O*+�2�K�K<��I&*�?G�E��z7�e�s���@�k27�6l`�J%z�X�s��HS�Ċ.Q�����[nCv���k��R�LU��Dđu>�T�ϗ�	��P����ȱ+v|�皏N�d$�{�1?��<LY�H�[���]��$��a�3}�b��2�P�~=B��>fT�j��5��<A�����3c��T��&�6�rD����>����]"��Ƌ��d���\=9���A�.�)Њ}MN�4��l�Pi& z McYE`t�"�g�v2�,s�|W�`�p�Q~P�N�֜D�{�^(�Om��~�l��x��nl���E�M�T��N��V<5���
#g�O'�R�a*Ƈ�|��Y�a:���<��9���)bm$���0~�j�;Ǩ���W(�M�E6�RF�"Ϳgq |�����X�$O��R|!f��kKV���' P��%Q�bƚ��[<C���Go��;�39{�~h�ݤh�Q�.�E�<v���s��Fc���"�٬_��GFЫ`}JX�	xQ~�%���Mڧ�}��	�sO*�[�t���#:9�V�����aD�l-���&Z�uq'o�\� �Y��`
��$=��ËHB���"����Y�(�y�\ʽ����?��ړ��C�>��$��˴1��>�u���<�/#A������bA2j�3nK�htU�(�Rdϑ�]1�yˆE�/�<x�z�c$ﭻ2^D�r��	�d�#M�.En`mr��b՜s��LSdQ�ـי�v��2ڒ`�Z)�����w��m�P���jNへ��V����BI ���K�
�oDI��[W}G���v��0�5&l���ggg^���"�{*@ֆ}�5ט������:4��_yMH0�e�9o�틎���uWr��3S-6����cE3��4�"}?�Y��	��t�.6���	Ǥ��|�ƴ �1�ʘ\��^K��J�Dѷ?��";�%q+�Ѳ`EH�����-��pq߸�T�2
�ǅ�j�G�$�`��ץ��ɲ*�"�-i̻#�^������2�c<�H1.(t�XJ���O&cz���ϲS#_t�@y�wX�qpؘ���	�7��������L=_�6Ʒ����@� ��`K���Vh�{ T��P���1RT�Wbw���z�q�T��n�W��?i�Dw�ql@�`�.�C�s�*��T��S0><F�ճ�絠�)ݸ"�p鲤��V�W��2�o���U���4��{�1���.|-�z�ǔ[��T{��� �a��m�7q�dӣ
{����!4�r|K����[t�V�P�Ay�B��EgOs��|�3��z�C��i�'��8 ���W���-Lw��Kn��Z#�V\���	ا�����R?c��R��/�υ��T��PU�u��ꮬ��|�f)^�Ȋ[�(cB�O���
�m\��3Mgg���fI5��}�{�WN	��M_O(=6��Ջ�:W��@��٭o�R��oR���d��`���Օ��]w_�V�ǫ�~���7ECF���[lbq7~��] ����O�N��a&l��W��I�2��`V�%�9 =(]5S�'�K��iY��ΤԎ�?k�4��X�	W����:&�2^a:���H��3�?�} *�(&���h������4>�&���z��>j�t�������B�iG毵�rBX�ݝ�L_��A�M��Td525*y�.�7=f�n'��j&�p� �'���[�%�_o�\��L�}KK׆����A|V�o��xð٫R��kɹ�
����4�)ɤ}��E�.f���9��p��:��,����R���M��u��xZ��xZ�z�N����/'���+�st���vS��qtĝ��g���`�q��(�ɫ2�,���\>��I�4o~j��r��(���V���&��"���N�,����/{>?&cJJZC��&R��3�$��g>���	���KHR��G�]�:ɂE2�ۙ�.|���7��86%�yw�
{�A���Q۝��5�bѷ�����S�~Ri|�v��c�#`W����>޺r��xK��!1t�	}��)V�|�d��*�����s��V;�?3�\,��IZ��_`n9�c,��-V�| �E7��J���K���Q:�cR�rHB˻��4��T�����?��D����6y�ܔ6��OL�T#
0�c�1ݚ� �5�Q�9�\��|�vv�?p%tl0���o�g�Þ�UH��v'�J���)WO�O��z����/��ou�'^��l=����[�eD����X�W��x ���|�fW��q���X�x�c�"��P�
���͉J��~���§�-2�5���Dj@6k�[��Q�[�6MN��sϒ���^��/�~�Lq);	Ʉ�`Q�/���]�8QeZ����OW�y[�ə�4\M�DW�����B�f���񭱈��D��y|���6��T�y0�A�!�P��d���˺>��V�[5�P<�p�_+��k�x̆CI����ڽ�(߰�:-n��DZeu~<�0r��1˝*�) ?�*���L��EM�گ.	q�_�VҾb�4����'
rVo�3Y��u�;ką?(����Mcͯh�pe��3�g]��K����ZW�c��<�a]X�AOB�ى�3$F~K��.�[����ꁽ+�aܶp����c�ҟ�$'A乨p�uM@��K%��m牪i:��_�I��؅����y� Ɯ<�
�8�mQ�+�I�7�]D��[�x����N�
n��3Gf6�n�W���_�!�{�_�T@MEI����X���T�������e7�zp��hOH����5=��d�����;��fo>��hO��@m�����] i��j�W.6�r_�H��,��r%`���ܷK�	������Kp900�����Ѫ�F�J��^���e��w�* ���e��x��&��_�ݒ�m�P:�L�;�=pZf<�r[9�I�g����[�U�?o9�m	9�e��O��U��*%e�����	_�Mp	�A���8���]�ѻa6/�%����놆y4n<e��v.Ud��[s[�"��MNb�s��=C�P\�5t������,��,r�C���[)/�>��N��0UЈwO�8xI��_i���?R�n�sx�E|��pxO�׀�_l{�Ȗi����������1
��e��th�[z-Q��M_7î�%hk�"ۆt�y������I���Ǘ��n�"��^��l'�p͗E�O��8�]��>���g��;��\�W��fT��xAL�!VsL�>������\�E���۴RwO鎃��Z��*]���\G�o�����9\�V_�������@Gf��6s����@7 Ґ�d'O_��+�1�Z��>�om=��y� �y �)=�W�rڍB睊+4��u ��Ig�`iĘȄd�	ۧ]fV���j2nu�
1@+s��n�ETg��1s*���v$>�~�s%S�M{���{�
ʙWY�v�1��Yt�7�q ��j�1�W������8��n��P �^��H��)���V�S��fc|o��g� +l��1/kt��x���y�7�,r�|`���sK'�u�(C�'��G�&zq��P�K;��N��E�Hr��t�<����m��ÿ��E��28�Q��q�B�;k��t��~'b*�`��``���aK����G�=��ҖڈC�J[����t�~��N�`;G�￮�䪚���G�w�����M�&�k%T��~AM�����>�!<�>�>�dD�=(�����tI�!vA��#w�VI��:n���VJ�Tm��	;->mm̓�W|6 D%��_̎*��4b�)����^R�0��SյTZ�� ��LQr����ߕײ���uZ�w]D�F�^����'�X��a<M�*��$�2?��4gy;Pm1�Э������)"���IT��/��0�M/���)�xe���v�����W�e� �)��5Aڦߗ�["��.[�=�i�O��Z���3�(f3|�r��1�����x�<�`-~ j
�t�b.|)��3��:y�*�haE����h��h��ס΋�� ��W�SC:�Sm�*���V-ah��L�?����|�N� ��m)�Y|�P�����#��f$�z�Iw���&6�ԗ70d
Ȇ4���uj�Z1�Q�_���:����?������0E�ƚRO�T�6e{��z׎J{H�l9��3���,@�.��m�A+H~�$c��=D�[����K w?���kg���3�Ǭ��&�;�9�9�u����]~��R�+vEO'7ʞj�T`���3�e�\_���iA�h*�S�r��B�[;6$	|,kĤ�FS�Ԫ��N�Ѹ�g��y��Mɨ$� ��bC5g�9����ݢ��UT��.r�q��*�i ��Ɂ�����UC��g�k-�n�?���5
�=L2k����������䄁�3{c�#NG�k��W�׮WW�H�Ml_���+@��1R�2�3��tpnY|�U���J��_��	/�tuӖ��il/W�h� K�ΧO��])�I`'zKS��Y���@����$�q��_=y��ڈױC��%�yT-��:�t/��?C���	�b�$da�H���<j1n7�]���tx��H���{j�v�~��KRr��.�������R葳4�|�=h���� �jA�Mâ<T.���������}����M�N��D�x�#�������2�[��^G��{��فC�d��U��[�ρئ��b�g�g_Qсf���8�;z{[�����*)rS��"x����{!�����%F�����r�L�	U�,	Ċ&���2���ހ���QU���O�;�� /�$j!�m�!�^���T�F��axM��|�l�i]#�47�X5�x�xK1P��X'���K%m��	h?�g�"'��"�%����[G��[�Ǚ�S/>v�Xۜw�K�G\�x��������SQXW��}�Kx�o��~���|%����-�(�,U-����0�`�C7�fG�.A:𔰙�C�g��96�G|e(�e|�|�mȿ��)�Y2��.IF�L9���������[��Az���-���W��2s�P�Z������x<[��;[�|�a���mF�L����i%�wd>�l���� }0�!���
��Sw� �o�ݏ]�_� a>Qo�\Q�1�������W���ạ�@	h�!吞�k�,���Ż����n��7�DU�?c2�侷�8����ĆˋI8�����QlP�$��㥆�zd���r�ְ�Κ�+OrRmJ~,7C�j�������}���>�����c��� �d76"v�
��=w���!eQ`��╼��~�E�.��S�c=�L�^#�$�MR�.}�h�ً&�Mh�	��,�+��(M8����^2�!�� ��Ψ���}�[����)o]!���&�$����@��祎�ꄵS�Y�鏈g�ڿ�@A��ߪ���Q���g�7}��S)y�t�Ґ�-d�}��p�OoI'�̳>:l���`��6�����ug�c_�v�Ӽ�u��oo�>��eg��F�_6�G�Eͣa�Z�9�7��	����O�ҧS�+��1COjѩi�V
�BʊΒ�f�u�Nfr}64��{_���nKe�R4�8��.��i$!��t������b��q�)[�4#�U�3�d�e��]�t5*����� Yd��A@�$}ҁ}�a��ΏS}.d�u;<bJ��u9�[C�? �U�aU`�K�����w��'��������p��~��C�����)l���K��P�WJ�L�-gn��Tk�[��T���mj�����h�!�ITŀ����&7d��Y<�����j�۪[ ?s��7lv���ء�zA�p�N9��`օ�%�[&p3�鄮�}D���MM�ֹ��9���d͢5�T���%N,��"�.�>3<�%'�"h y�&w����eb�� U�S��/��� �� Մt&>�K4�qƏ����a:r�R@DJ�����:��3F��]z�̀���W�`�����}m78�/�АA2�P15P5vA�>(�߄0Ɗ���?s��I�d���0���ҳ��L�� d�ܟ�N�v��_�����Nʳ
3�(��ө�ҝT3�x97���M!E��ӅѐL*�aS&�4��ᔪ��F|�$�J��i6�nn��X�M�u�ݠ�J9>Gfp�|<��ϙ�)�@�[�	��w�'B�Z�	鿞wX�{oF���k��c�r��ݯ��#�n��ɧꋱ_!�����H�cO�;G�w :}�T����i��x��>w��EgL���gT����X�vi�B�,��4
i.��#�~�Z�-7���hs�/�m'�z�œ7o�L������.L��]�l����ڑN��`�v�� m�Wԧ[�$Zc:��w��b�1Q�&����ʸ�h�c/� ����T,(��)�z'7^w����yg��D]�K��|�|p{wE!��E��lC��T9)�r��eƐn��3vnOQ��Z�d3J��x��qc�W��j����wu�?���M��.����[����(v��)G����S���)C�IO��p�i�;"wZ<w������'��!��ۻ��z��o&dӹ�*��ȳ`r}�ٹOk^�6�K׀כ!�Fa��P�̬�����d�n�@m����|���\�<���"y��	��ot[6��R-��Lc(����S��Z�B��%#8h��DnO4�5�t����hB��3��
Q��R8��b4|�e�W��a�jR��n�����&���`�\���Z(���iM�����g6�(�H?���u�ʜ�皪9�\�42�F%.r�"I	Z��?s\r����a��m�c�[7�r�U1�"z�*��� ,����*�� C]����o�P����0l�M�����xĨ�hX�	;���·��H�,R�(�1�:��s�?�xF�Z�CMň��^���G$��	��<c�(�U�=�*�E��;Ǽq�֕�ss0u�Rʼ��3���y�ʍv���Ɖ8U���P�B&�2"�������!�'�lRbڢ�.bsQ����?�H��q���H.��d��m�^Y"d��4Ղ��0&� vIT�rV�~�#T�W�*����=�?�|џp�WrrX$���'j��tW��`���y&�K�����0��ڠ�t��}#�"����`��+���k��Xu���Yk�TI�b
yPg/��6U�q�5 F�o���<�9���(~�g���@
��#LW���m�5��hjT�_�&�oA>D���`��y�I9JH@��=ښ@��>;�X�I�V�a�!:�2���)�@���:H�x2�2�Q�����y�粶�t��='����c���PJ}�Ő[Z��Y�uH� �8�p(W�ӧ���I5���0([t�v�K��U-�Ht��$6)�S��r3��e��x�i{�١�FS��xAn@�dm꛿`C��U��;<� ����~��D��z��0M_�
������彡<t�Gݰ	�6�]YH���o^�)XG�E���$0Q���3^�?�.�ս��7.`�� ����q�]E���1�K��8cU*
E`eFZ/��qcΘ��	gY쁲��S�K�Ǎ�Xy�����6�u�YHV�q[A������.�a^�zS0ҁ<�e������l�{���.������ 7Ԑ�y�,��ȇ�4�[�NfdY�#5� dV����^H�q�Uh�7����"�^p�Tz����;&�7�ʂ��_��l�oC���B]T�r��#��?i�*4���Lg\kCO�ƍ0�3X4)8:�\�_�z�Yn�N4n�)���O��Ey��.>F]����G΋�MQi����`ˆ��ӆ��K�[%3{���#�[��A��^B��Smw��|����y)x����=��Y��v64X+���Vġ*�+O��4"���0�V�J%Js���1ƻ�c��-G��`
�f�k�^��� ooY��X�㺓B�vE�Z wFݽjN�d��`sY<������ˠv�\3��m���p����obwۗ6�B�����muŊ�x�)���{�FZ�e�|��>��h���1�A�[Y��Op���=M5 w�	1t2UD�;��.N0�Y�8#��'�;#*=�>�iR���R������X-��bz�ߝC���r�O|$JӖ���8���[x��8�������^�]��q+��(���G�=B�z8�e(Jxo4a@&O���S&���,R�����'Dnz�Hs�H)sM��+��*�U�"4���'�I3�|����;��Ϻ�\"�����>���ס��Dn���;DELT?������a�|�XT�����X�r94D���Q^���(�\A��Eq�}Y���*M?�rV��NM<`w�ޫ����{.����Y�2!���)����9�@QQ(���3�X�(���{��Ī@x[��ޅm+����_b-���q���FHL���0ޚ6�E��ڪ�3�t@�Ղ1F�k*��g�׹늧#,��|�$iU���Эj(xu����`usM��le���|�<��P�$�N�˪��y���\@ui�1KZZW��WK�E��U�=�'O�4;�H�0>��V�t8��S�I~d��iF�K(2ҫQ���a1���.���3AbK��u��n&��#Dм��J� �����2���(Q�{�#���޶�LSOh��ጂ�Nگ2}��!��:4��N�LӟU�~����ژ ��G��@o��х7WT:*�����$�z�e���k��SM�^zd���$��`���	��|h�'��a��Sg��I�#w4Q�A�|e�N��ֵ����>���g�hN���<����A=�ݔ�z�t�	�n����
�O+�g���t$X�f�&Bt@8�Rblw�#V�(M=lL>��@9j��>�5Z��H�ϯ��̲} �M]I��V#�V�$\4K�J���3��W���/�ց=� ��f��Qi4��L��T)����鵄0�\���dպ�m�A+�Y)7B�}Ɖ/#��Л�w��}��h���r%D)F�.���v�n��]�X��p��[q�Z��l(5��8Y%��\o�+&>=2�3u@ u���2༬����\](wᦜ�U��i�IR/\�IZQ0~-�A¡^��ʟ�h�un��7��NG�$��aB:}��o�['ֻ�nG���iT��$�0W�;)D���ݠt��ˊ6��'�2��p�SL��vZ-{�ؠ�4j�2�{+�Z�?S�a��cF�j���(�7����:J��Z?�)PmC��4��a��@�t�ǧ��_tM��Ѹ����Vi���(� 8qV(�a�B�1�������%�K���3V�v� �j��TS�dƬ�k���*��-vm�cg�����!�*7�%=v�]�k/�7���1��D��JX�2:��,�	r�p�Ts�5,F�JW��6�cy܅�u��Uz���7Ӷb��J����kT��}���pC�V �����ZV�z�ٖ�����ufM� |�Ӹ:ozF�[���-�)w��ez$=0B6ʨV%��p�ڏȯ��j��I4��&K�q51��{*�ԥ�����<�M(Ak�R�!L3��.���B�PCr�6+&�E�~9B,]s�B��\]�P��G.���]��Ji~�`>�u�O�8!7p=@I�"�&�8&¸�������U���g�xȴg¦\)t�G��1�����~ѳ�'��`Ä��ע4lJ��X�ԛ!�����)��U�-)o^�Z�I4&�	�B�j�C��cR��rz��J�X�_��%NS�
��cY!}�n����D2i�6�ۦ�%C|�6b\������Mi��L��ѷ��r�[̟�ec��^���Nj$��V7��s�zM����Q涻�.
n6w�0?5,2�s<Uf4���W�in\�7��S������ekS�6���y ��x>��aݬ���bQ�Dc���������̍�'CHڜ�Kg뺩9�TĞ�ӿ^ŉ[��Ɲ*�5E�!?�@ܳx/�(��9M���_Z͙r�oҪ�'��AZ��x��U9�Nox�y�v���ڞ*���Z����R�gV�&���^gq�7�<п�yhj����(.��KP^���lK�_�W?Mr�5
&�G�]K��x��0��n���S�l^��Eb�ﲮYv�60{��F���Ĩ.�N"����9�~+]'�w?yHsK|vg3[x"�Ee����	�B�4�s��Վ�Ĝ�yڈ�'p͢eȳ�����)��E���JA���ѝ�幍�z��',Ųh�ڪzd4��Ɇ�ӈ�
E��L��AB�n3R�uV����olm_���=��P��.�~��� N[joi~[�=��o����YB&��1�����)�
-y�E������jW/�Q�a�2*�0�O�=ɜ2=��;/�>\8�K|��ߟ_��J˵�h�Ư�LLl�Q2�T��Tf��?%3cc��p҇�E7� 
���=?@��	p'Q�M(�7�Ɗ�^Ah;B$$����^^M�w��xog�kվ���f[<�k!��������]���K�H�ԗ��^����X��<�^cE��=�qPj�3zSj�5~Z��h-��� R_Ie�ܵ����C���C�`A�+#�柨Z�9w��Wr̜&H�?aǐ���$�ٺ�E\;THOˊc�/9�|��?��~aK���1�p�BK����s����A0l�X�K��E��e_4S��� ��$�0�%�\R�o5F�y�����P�;{p���E
���T�Z�7�����>UC��F��Z���$���i�91�ɬ�a�uf۲��&�r�Mj,#
f��M z��*0 �Jj����k:��,{�����L��(帄n�L�AY�6�+�����mU9�"��$���"R ;p�D�ʣ�_�`��
!s���/�b?8��	�8���T���ToC���@�7YY�~qD��R�+F�����M��k�ީ����L�c*��v͵�j���kN| 3�.���=_F, LN��o�pb]�tT�tR](�sa����Go[�uA���k�-�>��s��X���QFd�=�(�̈�^{�St�3m�7ҹ�M
67�z�B
,�I�����u?�w_�n���I+#��ڐ�;�hIc�'E`��Z��tW�n�����{@�����Kjөj2Jس������A��Ȫ��f+�rte�����vD(�l�O�������ܰ����7	�'�Y�?�[�]���&��{�a.[gg7v;V�,�Od2g�������B]	ɬuE>�]��m�@2�:A8��"��Pܻ�|��Fj���cЊh��J�x�՛v+��$ �<NKtģ��D<f�97s@�K�N�W�e��T����Cf�P|���lH3\:`Oa�t�R��3���d���)*I��,z:w�f(�(dc�ڞ[�d�k�򭵲$I�v�>^s�XI��nz�3%����؏����?j�q(�%}����}k�����{� ���I�AeA����y�T��֘Ϗi�����B�~�����X��ҽy톯��u�U�����7����dx��A�� �����1D��kYU�S��N��\?�A��n��>,��P�O�MUִV���=�cXʮYT�Ӛ䇉�׃Z�3��z�~�&~JK�>�d������	H���M��$ �<�j���<������B��ּ��P7�����I�42
&i��2Tu�����pO������fT9j�t�S�<_��r��RP�D��n���s��
j�9l�ͣ�N�A�������Z吣Q��G�:㜺�T���`ȯ��2^��3u����h�������Y+�[${��Ӧ.htbt���F{N������(s��D`s��,�\~%��ʙ]�**n���<�>�J~>���@�`���In�N�qG9$���B�H&�&5�Z51B���O����>w�'.&��IrW&�E��ڴ�l"ZC=�*���	��]a<�pE$h0�$\����D7��9#��(�/�,ho��R��Go�E�?�<��~���|be���i���/q��r��B&�r_�6ou�ݓ�A��q�����%-Ԝ���j��Wt�	�� ^�(���垤M��&��?��)�Ȑ�rt�}�3�w��dA���b`�:~������f�*'�
���R��t�Ha4���V��i�[U�E6}
��x�G��.��*�����(\�y��V��Y'��������I:�}E�0A��J�2���Cf�JUn�V�����S��vS�vn�OI�(f5�OG}�,P�9�@gm�

�-rDuY�2�"�5ٌ���Ee��Fz[��0H 8���Ǔ��z�U�{�}��S{�D>/E��Z\�Y�[�A�9,޶�S|�"���k���{f�`��e�5�G�=��ȯ���d^�}@"f�>�J`/�}��Z�{ܞ���0hz�C\�2�j����~��A���%'����w��.�+�r��u@�Dc��#�1`Ɗ�M��븍��o���Ͻ�c
�lG�	T ��/:��ㄘ����W���I�*�=�T�L3/�Z��Q�����zFrߴ�R�@�V3�!���-������7Ԃs�N6�V?�U��k�S?�4��njcA+P�WJ�yz��d���R$��lĸvv-�c�p�A2�xu���Xt���iʳΕQ��L3ؤX�q�Ɋ�A)�IR��9�x�&w����9l�o�S�n�W���#fl��!9�)�9%�C����uNxH����qx�:�&+�"5�cKkXx�6U-u��G,�uC#;j�_07�B��m&l�$V�x���
��/_	Ʒ֧g�UO����c<��:#0K���}��4����I��M1�]f*���1x7�]Q6k���G��3�b��I�R:�.W���btx��5��#ON�J���� �x��N���'Cw���*[~���l�t�.]i�t��_I�{��g1T�-g��WB8��3,7��ye�E�p#��6jL��x
��;)�4=�X�g*�F�_�S�P|�6�5�=��x�72�2����{��Q8Mfm���xW�l�����s�Xz<��8I���d���n�,��oSҌ_ͅ�nbK)�=l0b�;�(-��ik�÷->}n+B�m�ᇩ/~u���{�������_�����U.�����G�:&b�Ǿ���\=�אָ|�B��ߗB�T���)ɸ�}��|C[,����a�EO�+%����NC� �%��y��:*Q؇�/��jZ��L��b�����ꉹ��~̕�KL���^A�Wbm#h����g�� �[�YA�Ӵ����L���@�l��pQ������T5�Y��}��mlT�h��l���Mm��ul�E:�ft8S ��	�u\�[�)���H"�,�ݵ�ԱW���Reو9�.@��J#�k�0+�y�����'����[��%"_S��옉)��$b: ���]m��7���ER��s����Z�Y��#q�e������~w`�"����j����yv0�X��H(����}P�Ԉzc�Eoş�����'6�OP/o�o	2�)X�Ql��xw޺��Ņޣ�(���LS�����8���2�gH��k�cIu�;�G�we�E����y����1����',T�,��7��ͷ��6s׏�}�йqOl��CenF��>pj�3��L��S�XMXOOP�?��⹈�"����)ͨ:�<MS��,P��S�u�j ��Cc�=�p�HD�_��ap��l�j� ![
���2��P%:�e\���9���>�z�NP?*Y�hu��Y�6�b!�ś]t����켱��Np�H�ƒ��n���8�U-&C��#;o��5�E�T�yĕv6�T�gř(�@|��R�;�`���F��m^d�R�ʹ��E�<ַ�M}�B_�T�����������g���B�T���3m��ǵ^q
�;�8؂��M�?Q&�h�QT��9���]3��H�Er?F�D[U�!#�L����۷��<�dn�Z��^Q�|�wPo쿳�}����፟Be��[5�6�4<���tH�<=Hc��6i�d��G/�f֎�x�"Qw/��e�m���[a������H�!�XS����A o�b�=�B�� ����q��?��W=�IA��G�/�r�ǭ�2��
'8ej?Q�6)�ҝ����5����'��+ԕZ d���/�e���T��V`F�OS� �rw����KW;}��7
��B���%P�=���"�.h������4�����&�R�A�.H����bb��!#n�i�l`Ҷv(&ed��7N�3�hϙv�wg����R�s�8Υ�>�Gz�Jv������S��LXn�"�K*M�cZv�3 ޒ<c�j�\f<lN%@e�k�M*[���L�+Ҙ��=�'�p��D��fn�������K�T�(m�{y���ݭ;���:�:���TLLs<�O�e�w��+.zo�!(���<�V7U��[�7sI�H򧓒�zBVw&E$F���.�����hN깏kQ�c-��jĠ{��mhv|�A��2�-f���$�2���`j���T�1tA�i�@?������)߁�,y���b�lN�&~��{d�����.#G��`|��Y�P�j���w|#X"�m^C&�pr�ՠt�I��Y�	�����z��Ԓ�SsqC��g+�Kc�r_�<��[�����55 �o~*��b,x��Y7�iQ ������&B��[S	��*:�"�8)�%æ�[�'� K��0�b+;��~�ձR%����Q-9G�7ǿ���R1�����ܺ��5�����~�.#"p=DCHg��ՖibB�%>�U���ծ�<���G$
�E���;��W�?�?_��ظ���E�;-��1�DLy��rC0nX����.5Ֆ��5s��0^�J*ފ��%�)��5xn��xS�����^|p8f��v�M�G%�8yX���B�D�.��_s�$����A�[bo�g�V��<id���O�v����.��U�;0���!:).��͌\!�Y*�^�ǯ#3]��j��K�n{�@�_��B��thAo�~��^G�ЮNOg�{t����$�a�\�'Ar��gia��~�+�����3]Wv��0�E����ԝ�×-eL/5E�(lI��j"�W[~��pM��q��O�S�EV�A�Nd��w�:�l�z�������?���4 ����tωa�M%��TSق:7c?��`��<����̀dbm��|$�>�ր&�;b	3��w`�o�����fٸ�Yp�����N-k�b�h���Ы�W�[�fͪ�W�J����Y�(g�eEB,q��J��	D%GkB&V�| ��e�j�wU=Nڄ؋ ⶱ�_�j=�Ge����<��F�k��</�˅mee�v~/WE�-;f��	��@�0�5�[D
�g����s�a���1N�O-}��<���F'EPjǣ�����t�l�ok��dvT	���Rn�yߞ;���r�r�E� �`������Nhb5�!����k�U�n�����[@��3��ڵ���$�Ʊ\��;��	�grb4CJ��z���"��O ;���WH��ED*�Eav�!@N�
�5��q�O�NEhݺ!��ˇ8%�A���3��'d�3Z�b�鈜l��T��n4��c`F��VTLS�cq���W,�s�����P��n���e#�'b��G�@�%��uO���H&���kJ���;`��9r���t;JS����#�y=��a#����+�һ_�F���C]{8�ғǧI�)��6t��o�y�1a��U��Ϙ-񻑽bc�d')��L)�9�:w�}�2YW"�F��W�g�ܽ����C�:G�F���8����p�)X%w�x�,-���&ƭ��|pe�e�����Xr+3�R�,p2��g_��;r��<�o=m��6�� +6�����YXi�9G���*]#ފ�v*Ydar�0I�X�"����O�ǘs��oӡOb�h*�ց�Lpt�{��n#�t�K���� �Ew��K]�n���].���X4����0��q�i�

+ҟ��4l��d3�229���<�G[�a17�NsZ;���o;w��~��$/K�:��Z3���4A����&���'�_�λ��Ğ�Lވ���a��A4�h���w�[�oz��ĄwO$�	Ҏ�#7z'�hd��'1�n8�������݇q�W�I'3f��
0l=����L��ڡ�N����!��ձ6��_��\���|�aq���H�*Od��Em#��V�����W���Ao_>�A/X�� )�f}�F～�ݪ�������>6/��w�!�O�A�����dƿ4mݎQ�Ae-G.�2z~Z�N`��o�B}&��*xd�t��b!�DP�l��/�NHlG:�h��hD�OZU�]f���p�JG$x��v�Gfn�91��g�s�~�',� �׉�g5RR�$z]�U���E����8X�[;hQ~`���+"B���A	.v��
4(=��GJ;�jK_-��0���#aX�� �l���
��H,�Ĉ�h��}du�}{��78�����7>���<��8X�'
�#71����Ldi�z��w@� 
X�$�ܬ�,�2�縚������v���� +���p·�*��A�:�#X�PMo'.A+���|W�:�V��u\P�tI�,TÅA��b]
�����}w���PhUf��db�j�p,���{�!{�2�G�>~�-�'�b(���lM���U���/]��c�{���]D�:��}��T���ky0�9,-����o�[��uE�3ش���g�!��{���0,mk�o�ȬO���V���/��� o5}x#S/A?M��:<֞^����Vlߍ�����8>���j��J����pE�]��n����F[���<a��92�����C��[��Db�B�gy�Z�w��N]�w<�"�ֽ�/7�)��K��Iy�g��J=ɬ7:�X�!W�j�C����9�+��Jo���H�j��t��nOQە�n�P2|��{#1�87�.���}x��3s�~U��
��n�����G��J�>>�OE��V:4�bߏ�ĮB���9���L�]ʏӄ0�[Js���X(�D	?�a4^�q�#���,��^�ݙ�<S����5���$�ޞ��rd�ub Т�
tBԈ�|� �����������ܷ�V����.ȃ&�šА��1^Kx���G*��<lP��$q�Ks�<*��cRt�#�s(����yj�P°S�^x�9�U���[��%3�[���X�0/����2�8L�͈/�"�X���)[]u2m�G�
D4�F���V�<���6��,I���?�F�EB
�o��.���P:<���L��-��P���ύ{V$�� ����0��׭��Z9��.l����V+�hA�i�	��CX�Kb�w�nʨڀԴ���2�Q�fFbx��ЍO<�>0wσ&�r.&�_�vq9_��*���F\1��<�B�(���&=U]<�m���AB�j���S�Fzg��ɀ�jt�|&���)�2]`ϳ,�V�q78�~J�G�N��q�.�1��f� ��!C���z�u�U��|��z�FN�P�|��!<���m�����Ս��N:SNO�t>'L�}w��S:.> 
�C�vt/���\q��;\A�6��+�[���q��m��	p'��P�J��������A�ހ�Nm�r;$*�o*NM��s
x9�  �f��O�+՘�Ҟ�8#�H�m'��g����k8�d�&��=O���%4��E,pInv6_��?�n���K�ږ�j��=�w�0��x�w��1,���ps�4Q0�"������#4�K���"����H��-�:�X��u�>l_��(Ƽ$��
a��D��4��ԣ�	B�����L;���Ml'⡐�"A��ҒRx3�!�?�^���3�B<i�N�M��ƮUqx���Hsj��~}eZo�G4�\��
Þ�?3�����V�}5H��U�T�'��cMY�R���]'�����M�7TO�𭳸a*� NG�Mw� �z���B���&�5�e��D�=�"Ad���ծ0Gړ��+}�P�~�!�:�^Cߤǂ;
� bg9�V'���K^���-5�U��!!���?�s���L�G��6�����#����-�����0��{(��'�Tw�kg�M'ev|�x��WƩE��.�}�%���\� �O|8�~���Q"�	JP�`G�vC���W�k�T�@�#�4u��C��T1��iXz�^W�-��ǰ��^��6��$�䄁"�x��e{\�E����|5�.��/��jԸ�8Jyv8�1{Xꮫ!i��:�0\������B6�s%��������B�j޿哘�e��	��Z�|<?uqQ;Q$O׮+��{ۀ������e	�B6�1T�޹�5�RI��s����irU�+V�z��f�s�A���v>4Ty�F��Qjw��C�iV=9D�ɑ�e�,�����4��(�WA�4�����F�י/:��4q�\;N�]�F^������pc�+�`b�巸?W�p֜���X��_�=;��5Y\c=��EOk/8�R�N����V����/�0DK'�%��W��S�u��Nb�>�ꐍ��������5�$�[x�A������ؗ�hlaJEp��7"��-̲G��.}��7Mp<��E�4������6搦%zN����7_�9g�� e�ڸvቹ��Jn��Nsdɯ5�M�t�KFF9��?�E1��I�?����i���+�����a�0����(�p-}�ފ,s�?���I�l��,�+I�j�v!v�C�b��	�,E�g�\�C��T�k/�ަw���.�ȣ3�l���7��)�΁�`7q!�+�V�g�Rj���QI�)�������\�Y+0�O@^�T�����Nu�_�8�98�U�a^p��E���B��������`���*-���/�``�&���
�6��4!�]9[�-,(":��m���N��5ɱ܋o����������<恜mlOZ��HG���ƗRy��JT��"���ckGB�}�=�)� p���O�V
L��Ka�eϿ[������p���U,E%+���8���yj3R�[΄sk1὘��#|�����i*����s�!+��JI����?M�j&��N��7���5=�����R�cW��qRNM4���RD[����Չ�w�JҔ�i��A��6RZ��)p�������J�ɥ���5�\�
�A+g],`_�:]H�+p3�� ô?
*��*�㋠�1��c�ͮ�"f�E/�T��{��R.�h�*�}g�1�.ɋ{!�%�4Xϻ���9�3H�FJ��\���?��� �Z��3 �d�Y�/�ysS�v�� +���7�f�%���aaRD�:��a�V�5����$��f�z��q�ȺW�͜N�aw���?������7�X@ݹK��V�Dy .��"�+�c)H,�0��Q�D�@|>s����>P�&5��>����y(0p@���������z&&߿#Aʼ"��0<C.q�f�ꍶ�����	%���7��+|�O�;-8<�^v=�M}����pH���/5���=iݴ�VCDY�V� �RV��MIyci�;�񟗏jK�5kC2�n�f��h�,�.��{]��|�yQV}�TQ\��~g��D�<|�I��U���Q+R90(��M:����@5��������CC~F�j\Z"��C�v�
����[s2�_�H�51'�j����"�ģ���|�T����au�S�([Z6h� ��<rPU  �=9譖53�����O�ܥ���y�_��XfU�ٵM�ˮ���͢��LC�|˵��M�]=�hF8(�O�rЩ�|��9p-�>�`��|�v0D���h���m�36x����4��+����6�9�؆��N<����1�1��7�H:D����?Q�����VT��d@sc@���~ΜFF��#N�� sbw�j�,)3��/�	�n�ݣZ�1}���	�5�	|��d����K�𮹷�?�z(�m�z�5�󄯶��Bg�T�^�@[�i�F���2�f�����n����I\v|PF.0��6���DI%��;١���=м<���I�����}�-�'��mc��v�Ycc�,d�k�fK���6���u��6O��B�T:�Q�n5�/(�˫_�fK���!]c�bX�E���##�F���Jy���5T}��J��uS o8��	��'�;�h#��?r܍��8f F�[Vn沰�E����ZgcBjdoIN�NkL��(�Б��"[�9'a�j�Z��	DR?ȱ��}��.��I���5�vom�]0f	;^��"^�k����:+#�c:�ڱQo�29���r4\��h�	�),�ϕ)��ɗ}D���t��'-�#,�%�T��0�Ɗ+z�����>�zK������=�����-�4�,gF��`@�N�����տʾ�խP{�sb�ej-bj��1�P�)�$qo���%�d
y�Q�t^� �]m�l���������7����<��9��ʪDE#���<;�	��+�Iw��~��w����PmEkG-�}Q�d�;����{# �+/����h�޾��g��
DhkC��
���gbɓ�ϰ�v����`�
.��8[�Yy�����X���������O
��J�{��3(�%�;�MNg��Yf�>�,��Vuď�u�"��ȍ�Y��G�#���9@q�M#��w���W�uok��G%��U��,R�h��xD����!��<�`�i����R+*?�}��'&7�}.�V���lr�w�}����q�
47w�Y�����$��9�G�{e?�����j��^�[�B��M�����^�cc�F�&3�qlV����B����"d��h"�)η~I�� �������o<�ap?X/�n�6�f���L�R4˥�Hm��R
��s�2 ���.��g��>�z=Ύ��ɨ�^�������#�����*��ۅ���K���P�:Me*n���?�؉(���N9ٍ{?�7^�y�RX,���B�o(�����9���1�،J�.+���V?�"��aVc�(��D��Kc�X[G����&�|��
4}b�4.5�n,�T
5���q�>� V�E?FyV�(���sNr�>W�w���D� �U�p��w����n��$ƺ����b��0{����0o}̤=_h��$g�(�y O�ݞ�\\6\O9L��ߝ�S�xI)B���on� ��L~ۅ���P�!�!}Sw�W&����K�!�;����,��0�SFAό�n��RF��Z1����hc��QջglFU���[/�����ߨqgk���&��qQR���L���2z*~.�(%���C�e��]�Mqj&��dڻ*2p���po���D�Ps#pH3p��ښ�����ս��'�W��cE�@�?�L���6��z�g�L���Qh�`'�#K����w���ٵB��nj	"��v�͜�@픾%5cJZ��u�w�2��X\�����|&����%���w�d�-S��/eܛjQ��N���g�	B�Uݞ/��$��]�����6
H?0���`%��=Ģ��v������ֳ�ܞ�.ߛk�r ��t�7���̶8jkVIXh�1�9��c&C����W���9��(��Y���PH8u§��N���:Ӯ����/Iq��G�|��������!��t`9�Bώ`���ܿ_ԋ"�*�V�����2k�ڙҧ�8�y��]'~Q�«�.ʈf�4Io�P���<�øUZ�%_��u���Â���e��~��U�/���Zm��L�?�s�˶�f�M��Z�T�� ����+�rĥ�Y��Hp:��7�I�U? x 4��s�b�R�^�N6 �~&h�c~�F�)��b�s'u�z�����T,��C�����''�(f�g�Au�� �T~��:�ϡ[j��~��I^���r��zQ{	���W��$�>|N��y�A$�w�}�4i�ђ�\,'�!0�S��&�����DC�7mq��̘}��}v�}4(��x�l�_��l����!��I�G�,P�������ڟ���>W+=}�'�l�s�SP�G������Ⱥl���%j����o���ڰ�~�q���peKF��/ʵcď���'bZIt��;�T�n�%p���Ns�Um`<�%�i��ݜ�z�6닗gQY�(�(�*�o�d%N><a�+��H����|,��yK��yZ橪Я𣖥��!��纎�ӆ��w2��d������.�͈D���
ěa��vTt�m� o�s%(�}z��;�L�t1�K�HB]-C�*jQ�7��=�ɩ�d���A\H@����Zׄݥ�I���j.��إ�������E�n/$�(/�F�%<��ޒ�0�8oYfmْ�#�+�2M,4���5}X��qZ踎�ڪ����H�a��\�|/�{��6�L9��N)�Ӫz����_�ư�Áp�*�=v��H�\tn�Շ?^N����Jw���>v�"��y�I;�evf�E孵�P5��gr��gɾ9���/a9@��T�g��b��F�"�.M�e@(k����kjW��<�P�7s+\���2��P�T�?���$;��m�Mn��dY>Zzd����8�L'��"ƑX ���ӣ�g�/����},Fđ�e�%́�E����!C��0�C3a�� �f;���H&��J��|�J��h�\X.��ɰ��#/��{֯���½��$m'0C8��vqd���tx�p⛢w�g�?��PXЙ@wĂ�ۑ<P�<�u|�Ui�?�U���G������\[���\v)L��_���V�zZj[�Ơ���͆<j7��9n�?��)=�t��L^/��}
�o��e�4o�/�^�L{g��X��"yu��|����\}T�<�[�QP7�l�++�"ֺB�2��A�Z,�n~���s��w��𲖅�ҫ�U��np;����Y��������T�(t��x-���t��`Q5�Ȼ'�8��p~��R}BN^t���Dꁘ��/	�F�h�k��݄�zn��w'FA�RIԌn[s=��!�����!�U"}ej�*ܹ��4��}Ul�^�]u2�&ӵ*�|��!,R��	�خTN[��3 �m�.���cN�����Ge��m��ے�q��a�% 摰`w�y��M ��[h�M�'�_���cI�:[`y���ӣ��H�3�ށ�����U��t0�� ���s�mC'O��O�3%b�87b{��6*��[���g�T/�M�!j�~F�����N���)Jɾ�u���s�~ߴ�� �eu��O	A,�N�S�JVtdKE�"��g_�c�o���[XZ��ˋN��VG��=�^*Y�QzY���4�Z�Yn��BA�'��~�E�0i+xq��w�b���k-�wuxp�XKe2��q�
�,�?��#'��P�RV������9�W�nR������	�-6!]�����{����+@���]��1s ��ta�@<j��=z�����XDDc�|R�Ձ��n�FaG�C��k�ZR�li���ڷ>#r��b��0U���4s��Q8�~)9؃�1s��s��d��,!5ZPUIr3�Z,D_<i0}=7�e[������HB<n��'�z#[�5/���&D�j�z�^�n��*��;j-iA������VtL+�qd�.�Bp�bܼ+KK�Ҽ*���[�B͕,�����Oµ�B'��g�g@��T�,�V��@�d����d����_�ՠ���잴
�����WcA8U|Cn}�`���w�Y��T��7��}�$�,��@�M����.y����7.��*=�u��m�.M���/�-K�Ǟ�|�v\����i]T�#^�X����e8RK�̋d�X� �Ql�@�h�k�e�|�w3����~�(�g��$6�>�Wv�K�hP�X�@y��ߖ���	���=D��:��
���
)�n������_jJ�&$f���!�OC�X2U XJ9��j���˕����2c�箮����"�!�����Lg�?��>W�[Q�I@y�h:'����Y�! �Z\w�����L�\h�m�H�Sa'��Zg�E{���U��9r����?w���Z�i'�q$i�Rc���Z�j񍩢{y�y*8�����Tm�$&h�+�Z�OB+�9ҹ���3Xv��NC��%6�4[�EPk�'�I�(�M�rK�_�+�iq�3�R�	{b$5��uk���a�
JIZq���K�.����s����/I��v��&���� �jp0��ս��J�^��eٯ1SL+��'�KT�Mp��S2p8^����Jh�������lt�Y�V��C��~Əd��6��/js�s���ΞvX-�������p�[M}o�g�G�uS��(���'��_��y���G�ݶ�]�1a�����>C`��ͧ��&�<���I�1l��Ȫ�fΡ-��GrJU���qM2C3̤��`C�~�v~X��i�n��E�ǌ�r~4��<S\�.T��/.��`�Y0�?R)"4����ލA땕�)~$�K�֩8Ч�J.�@�oR�>�IO9�(�[������]�봺�'$}����^����-�_����W���A�yaM�pqz�o�~m���Y��7��.��"r�.`s%�}�c��i�����ӧ�LK\��U}ttE�0��_�����Vvu�q��B�)X������c�h��m�>fcb�=3�͠�Z�R�厴s���|JZ��=�ڱf.x�b2j8V6��첂G[��F��Đ��y���y��F�k��w�YҊ����tl�4���Y����9�G#�.���?j+�S���g$1���f���P�<b�.:� v+�Æ��+ �LwE�C0�+ڵ�fM�{uW�����.s̾Q��J��R��V�ҙ�a.�
}�S�別�H��M�׽�>τ��ӖB¤�D�:"�_IX�x��)��J8�|�&�{���ޔ����;���nж�j6�F��E�uT�E���T�������i�S��ũ.Q�D�I!�b��cR�V%�I��Ւ�S$��Q��~v���n���lC�'�!sg�������c�[L�<����gXx�_�jӓ���צs���-���ӄ��7�5�����h��G:0� MS�F�*{b3�$/�3�}
6#��ٓ!ڄ��j���%�h	��H.U�9��RB�����B��ZRP��*�}����J�8�pܜ�-P�E��)6¬+�Ou�ɖ���-�-��'n��8���"��ɢ�_%�;~�g�͝8�!�����P!���.A���B��i�U�n,Ӫ<B�'��\K����h�R{V_
qiy�d�Eǚ���ga2��~�흮:H#`l�j0-� 	Dmi�ST7�2�xF���o*��
m�\�d��9�̂���ܹ~�X�ua`���|-�!l$�ꔺ>��F)S�O!���.����#��g����n)H<��-����mEm�7��ȴ�.4�6��ߠ�����iX�a���+w@W��*s<��ҿ4�b.u�Һ��I�/��^�����L�K��Y+"��zl�;�0`7���jQ�@���Q�v�*�/Z�u�2�7�[��Fe��.�m�Ȣ�=H��#�Z�i�T����!T�4qר���-S(�r�^q�PO�nͰ��j���:;�:��o;�bH��)�Fz;c�=��N����YS��ƈ�M�Oӽ��:����r����{�Eτ
G��>�Y��[g����\�g_�����9�<J%�䒨R�	#�W=��~���Z��0?��ԓ|
��H <I���ࣟlc�q��JaD���F$���[�k�l�z|�%(�mj�����<+�����ݸb�E�6<�C>�����-�;����|�zA��5Qzx�Y�
aw����&�� �#7Tc���P��9���

������v���F�G=Ol(���'��ʰf����c��Z�ϛ��gr��@���?}��S
#�Ey�I���<��w���[X�����e�O�<�W����)5�My��Pa!��`���oqk~���ڇ�>�4ӕ9��$+,��\H*Y7
Y�9�x�k��0���&E��DN"*�n� �6���zʼ�ymяFaꃎU^V}��t���I�mȲ�a$������! �{���1��@��6���g��xB��z7� _�֭���*}r֏�	�f
lQe.@ �ܜ�*A�O��3��ӏ�yy��5���
��2S����zׅi.K��Ԏ��G��w��?�]�y��RFAú�k"�1���\�n/�W����8*�$!�v޷����o�U<#�����+��h����=O��X-V�����Ȱ�B���O�fD�]F��)�kHBz}�g�T��W��>oP�M�I��ZV�ٝT��qkDEҠ�S��F4!�\�G��A��85�2_����7�t�n��Ԑ ]LޘDL�4mo]/��+.�y��R�L�b��&d-Eok��T���|���[�`)��xkːO�����z�ن��E���D��͛aS,����H'-�:Uw��_w�k�N��]�Z�-}�l��Dv�;����W��=5b#��9]Gˌ=W���*J1f���J��;.��9e����Z�R�4F;���W�EOC��*��#��u�N��2^���H�#��O:����X�1Qd��K���d$�C����Wfl��(�F��#:i�Q��Z=�f��o�ٻ��IP�w�5D��;4��W�<>V�R3#H�RZ����/�ѩ9�r�Uu�)lYu�UCs��O�����B��w�SM�sg�#�h�L�$�pTU��x���j�(���|{�0O}���$	��H��|R�ϰ��$|��75S��q��]zB��6G�Ҕ������ä���FnF�$,�B�d:������<է���{��ȗW����a��� /��{*1�P>d@a��kI�xU�ubSK�o���, *�2��hw=�D�k��|�M��D��Z��c�c�5H+:0网���I�R���If����'�w������hx��)���j������r ׷J"�������nR���I��՚`�#���c����)���T�q�Z�R=��a�`��x�yǮ��8��fo�-�1��?zEX?����/�;P���H��2,BM�
��P��hG�6KF�X�坍+��9γ0y��A�|��څc�A����Ges��%�뗋�2�/n� ��[]{?���9����VhK�"	�Ǹ5�����U�si1v��3x3�4�Z"�E��r\�!(��ܻ,4K��C�&��w����$�{�mP��'�Q�o�R�͠D�>�C����^�����İ��q����������JJ��#X#�^S"!�;>"7n��h���Q��w5���
Ü{�N�5l�63��vv-Z��
�{yX`$k�f:�P���1)���e�K'�bFXut(ķ/*��^c��U�3�%� z�y���C�|Z<���꽖5 @7@�JM-ל�ܰ/m/RB�BR�'{��Wl���n~$�°��A�h�k�H�^���eٹQק�d�	�Ki�8A@�R��
��sr� R�[�Ţ'�S}P[o��u��$r��6�v;�j���g��T�������~tv8T�*&�)������ eJ�R{N}�u�S�ìb�c${jx~�"�W�H�l2MLe%�w�B������C$�Ƒt���4�8)c�Z�-�dlj��a�>�U��*["lp�Ό�J�vG�*5�D�MЌ�`C��Ƞt�� Y����T���6��\���;�:���]��W��������qd���(7Z���F�dw(�yI�ދ.1տK����\����b�~�'�9Q��J��r�=��0'()�@ѩ����f4E�jX<ߎ��a�k�UB��㾩�uL=S�/d�"w-�����9��g%y�$�W�]43AC��N1�4d�u�C�J&Q���x-[�X�id�	9Bm��̔��샞2=N$`uQ�H�;n"��0��f��s����R�hL��y�.0w�4�}d�xd�w�U��@���9V�ڊPk�"[4�	��y��s���/���m��V�_�33��g��zMU7:.���+����M�|Y��
R�$p͉p�i��! r Yՙ�oa���nԔ}��$Ƴ�`-�����Ǳ��Cg#P����oF��l��TG�ח�D5隘�!�����IAm[R��4�!�n�) �+�ţ�f�./B��t�'Pm+��Q"��]v(ٱ���nF�<��ʉD3�?(����QF���[Ɛ�/V�<6,������^��b�&�cUb�;�?�w��>�H���>�[�Tp��"���O(@�;�k����7��]�-进e���
��<փ��j�2��CD#��'����%#z�w�;���Q0�	<;We:x���6B����(/9c�i�ΓDb�c� ��e+? ��v@�?�#�9��U�]�������$3=-JV���R$���b�R�~}s�U]�צ+�/��?�(�F%/<�]�E(�e�uR[�m"�8�-~l��a����I���t���}�ͣ? _y��6�LXPL��ɖ(���0o��Qж�no�oo���76�h9p����;)s�5C�)&w]iԾi?:������~��Yl7�8�M�`�`U!�Pp��x�6�b�s�*�_�J�	c�Q�����YM�Ж��	3M\�z�l��KĿ� �	#��U�����|BK<Vc���_ ̒�k)���<T%�o8�|��+{���`ݙ����Q�IҜqy8s^R��[�{^%���[8��4Y7y�c�>�[�ɒ(�$1�ί\�ϖ��9Hv�Qd��Šv��X���!�v���GM��h��`X��cd3��w�s�.�9�_y�!]�;G��eP�t���ם:Qmmɔ���l4ځ�@ہz/I&@
ߢ�1�4G��lCc-�k,��o�_�ܕ<ed�!���R��m ��v�Ɣ2q�װ��ԯ�S�p7��}z��� Dw��̢>�j����Iz�Vg��� �Rx�$L������J;�]X�%�K�2.�#x\�0��kИ�`��t�P�H�n���6����!�C�B�'a�Q���L��i�����W�bx��¤ꐉ�xXP%�ӹ2
��
��W�A��s��kg\��;�vC
�&��[�0}���[��:��_g=�A"�H�����m/p
QCUc�J�(Uia��
��@� 4B��Vb�U���!��=��{׎�E����\W�Y�����nF�x��;���Ǟ������(�C�9�#I�p4� z*K�~�zYO:��l<Psn�C����U��RymY�6!�,R�}pd�4�υ�q�(~q���u���-\a����ͻƨ�����#�`N�ǔH���Ƴ���2i��(y2���� -iX�q�������R�/ �$`�G�D!(��`N#���o[��RzM��_�,P3O�G�M�9f��I>��!f���i|�ʸu�a���W|�ҦB�� ��`�����ޞVJ�I��/Z����\�6�F�s�z�id�O
bi�y]3M+�0��q�&Y�ױ6@�V���$j\I>\Dڧy����n'�b3<6��L��Tx��,X�H%
�������mF���儒����Jj�Q�H�)cl���q�J U�C(��~��0�E�� ����[/��������w��g�/�蔱�d�
� M��^�s�N�\�_/*��7i�1�Q)����x׮N;F9W��4:{�Ɂ��s�о�7�r�lm/�y�G1$M��2�*;��U��a/��S��R �]�h�rZ˩<3_t�K"q�V��.�&t��#3�(�t�Z���׃/�[�B�D]{S��$����$����y��������w��e!���\T;��#��f}�N?�Ekd�16��ps��r+���&,�#\?�X^�w1���� G:�*sw;bj�S��u`�e���I>R�MR��?�F�r�5���J�a��Eߌ���[��͕�D��\�=��L)@��ä��-�}�&h3��f�7B �u.�%�@Q-I�uw�|^�[/I]^��>*ζ�%����}y y�m��ëB��H��VKVQ �z_�Ӻ��k%ώx���.�w�4wq���_Y"/^u�r8H���X=�'n.�����	�`z��@���AE��Y����<�j�$3Ӯ�@PIE2��Ywg-�;FY���U4ok���-����1�k��,�=��Ɣ�N*��d�sk�y~��8��՝�v
�&�����-S{p�9/l-Q�)�V㙘�:���L���;�335(v6�X;��-a�Y�tg��3��XE��qL�t� uSLZ I� $���� ��q���ɥ��W�������
����6?�r=nRNBT���B� �5�@+#�-2 �U-؛܁J����g���1@]�E����j���cZ��}H��"�.�cZ��9Z-_�[e�:O}�Q e�$���e�R�bLA�/��E(���%r���o��{�v��bÂ�c��8��}5_3"i�f���ƥ����BJc̭)U�u6�����Fp�C�e�8�<����)��ku�I���R�7�-N����4�N�,�W�(���j.�AV�R��򐌫���⫹ �I�jC�Y���tdŌ,onzӭ����#�,1� /�7�������[��С�Q�*�t�w j9b���eV�Yb��I�TZt�����$aCENS��I;�s������T�w�t�X8>�?����c���7�X���cߜ�Y�_�o�vlL��P<�w���N������'�6�e���T<�h����ݫA�8		h�p}��T_q���=^�j����}��x;�!R@F��H/�Ӷ�������	(�g�bՍ�Q��^$>E��?ܖ�X,#;�����4�}�5{Ӣ����Z�Ș�ٞ�EԈ��-)~8F�A���p������*Y��*�V�L�K�.
A��t�Q�x#�9�K�:� �i������˻�6��n���i��7�8�p�F��N�0�:g[����OWx�y�ok�9�]�ģޢKiF����X����a~H��d[*�0��� ���%&�f�^$� |��N)Nz�mQ=�r�Z�e�ܳ�����Q�T��HDת?.&�"*��������{��j�VڢCN(�w�d��-vf8 ����d�F����݄-��[x����B���n¾����(c�6|�K�� q����(p�3��OSO�{r�F<$vb�lYͳ�ӑ!�f�T�*�JܩZ�GG���z'<��Ia��k�Y`�Q��%F����I�
A�$e�z�`G�a��V�B ��R�~d���FY��l�;�/�@���*���}�C��X1�'A�^����pv>�AP�Ù��`�OOr���Ey��]�m���m=�g���l��3�#�I���*�n�9�Y�.�����n%*n��0[��Uy��TB?:���
oB����&��s#zyB�ſ��|oR�������?��?�����@�>�����vZ1��D��A��������K��H�|1{��f6��b��:��_Z5- x��]S9�T�jkf�\�1�vw�����Z�G^>T�n��i�k�zښ��O tj��R]����"Iz��  ���RW���}�i����?l������:�����8,}��)�Di�w���X;��!�r����w�]����P=�	~=�-���af:�7�}3`��0�u�>k�|N�r��������J�th��j�e�2:p���q>��a-�r��c�v�:0+����\V�y[�ߔ��J�Z��0!u�w�	���i���.�@��M/c�����8�.��$q�򅉦���g�v~��Y#@�����
+�6,��ԡ<��e�{��gj��`35.�n��k>��H{ԥv%�hm��'ْ����[���,��]>��e��3:�6m��vE�s��QTO�fs��g�9W(�oZo�ߍ�b.�Ĭ�{��8�Ť�|}��.�`�����-?s�Q�F|[���6cX�j�$�����D���͓�Z~��Xo���x�k]�	d���K<p:���F�a1|��Љn���:1j�����[��w�bJe���.�R�NNI��H�vv�-lIM�:$��t&�xֳׇm�2v�^�5��'�+:�(�P6Ո�'��2��~Jj>A�]((��e�k`V�c\Y�;B�t9�3�u��Q$�/E�L4�,�	�=�*���2��
n�D<�ݑ7��`�I��p�j�P��|�a0!o��{�/����-z����Ā{X�M�ځ$�3�e:��?�!�_��=��+��������a�{�&��j�a�a�e�1?CN8����M+h�	"Wt:P��ӀD\0]���:�h0�����!��hc�O.S]Jb�d�Va��bD��a�؍���Xe���l�क़����8��X|j�)@!?_��2_ԔnFUP����{��1�z	3�b�a��k���-�}1��-sS���US�%��+iu��H�h��P��.��'Oe��u��k�|�k�>3���W=}��7v��?���OUxs�)2Z�ޡ4�>/[jL���r������<����oI�9��1���xQ{C$��R����;'���}��%����>6���B�3�n�P�.��0S��]�%���M�������*�^l!&�1�,��ɰm�H�-22ϫ:(�����[�%Q;�si�Qy � r��� ��޼�Ś�Ե����F5�V����H�0cvUv,���Ä)zkk��V̊�ݵ�Q7h��S�U�ʬM�W��'#P��xyC.`�8�҅/c�x��{�Co��j���|틼��{s�뛚�+��,��d��Ug3�� z��e`{����q�<W���v�WϺ�w�B[����c�ϵ�KOت��0X�W+\���u+���C�3o)5������@h�=L!C8��H�=��z��	E��T�%���}d�	aDY��zG��?2�7���/%��i,�я�5�.�a�	�S� 9�?|dk�I�l��{=㧌=EG���5�{,���I�4z2}\����|p2����
��i7��<Pވ�+g��Z�?�l9zvN�� .�щpx�8Yź��1�����R:���h�РHId�MĴ��*�-�.�;�3M�y��ʠ_"�c/�?!�j�,������;��R�h��zE까�Da��j�-��� n1:r$���7��D��7\3B0
M�ٸ�nE�i��+�*�H�U�n_TF3�o*�{D>f`ض����9����K��6t�-��vzR��q��5}ai��" {�R������9�{�>M���)Io�Yi���a�$�5���$��D]�LV�A�#+ի��C� %<(&��QH�u��Cjkӕ}4{V�<��xg�H�̎����Gq�;AoT��$a#of;��#��~n����	��n���h�Oć�O�##��HE6���"=� �8�V�\|��̊7bYm��?j����s��^�s-��,��ZA�������V˅����o$.1^��%4�D6D�o 
��_]g�p�O<r�Q��ѷu��8'{�ݑ�p��!M�P�;Yה�r.��ɽ��[%IS��P�x�3-ɊCf�(6�dy!����`^hR��I`9؁�~�wQ1��B%�^�R��f���p�C� �X*סk�\�z�ñ�yOÌ�������
�1���Zl�������r\�\^�6�-�}���\K4YF������c?{қXD'��jip���%YYeL��%Ǒ���7��'�h��s��T��n�Y���R����l7�sz�?�>T2�^�{B�J��6�訂����dA-�8&z�+������50is�!�^���ŁI���H"�뵕�P����hk���9���.��QK��}�&5�'�,���s��gi��b�:�mu�"Jw�3��=�M��$r)^/�T�t�9�c(�廬 ``�&����C	*��TvJ�n�d�6X��`�:'
=�g�UU��f��<�������N,����AY�&uD��Q�OEI���Ƀg[��Cq-��O"�ܗ��v�ֶr�^�%�oX���	dKcAwvh�%Ѷ}����&Q�'�v��^p�e�-z ��a�f�R��o�8�G)u�,n�*D�����+�o�S�a����ۗ�u�_���'��_;��9<k.fge�樀@,��d�v�C�U����l����j0 ���#j�������^\B^θ�%S[����1$d�dpP�9�`��5<&1�Kg�CǬ0�*�9���݇��I{W����Nf)Z��`>�sy�W�b�Ǎ:�g+0Gå�t�$B�������������>�F�1;�8m���r�2}�c��ʭ �MC�`�0��!��Y�NF#��`��� L2�S:�m�0�
:�DGCـ�*�D�դdӊ��4P~�|�Q��O��5��^��UZ2/iLA��e&ōb�Ge�����jx4H�?TՂ�-̍_�L��=<�CKo?�YC]R��ØdBGLf��ts�WM����&��տ\c$��������$�I_��Ao�H�ާ�%�9��(ء{dL*����H��>ҹ�% &�c�q[�����D�Y�a�u���� �y�tcc񠵤4�n�"��������%��@E 79(@JIw�Ȓ���f��Xd(��	��u�F��N���	��ĺ�~��ƹ����A���2��J�p*�i�G���?�`���f ��V`W|�<^8����	�F��^A4�%���V�b�6I��X	���b*�ۧ��������oP����Jʱx:+<\�ܲ}te��ǨWN�*ꀪm�{3�+�XI��7gHMƀ�Fa^���_-�;@�U�\�j�m�l�+�T|�B�<xM�Ua�5ъ��7F�R6�o)�p/-��v��3�����BdYcBsBQ5Ni��&p�D��~S���*k��m��4��6�Y�k�R�4V��Jc�A�h�׬^�G��<b��
aE�����fד��[Y`0�ɼe��y����=UÎ"���%Y��߈vF䭸����ҿ�
P:�v�Bb{U�x8�Fv@����C�'���!m.U�xx���P�V.@���
� ���^7D��[�ˍ�
��N9�r��T|�p�U}�6��	�������E���vT��&;�yQ83�d&�[.:CB^�����C�iof���c��m4���m1�+�*�и�jp)ǡ��YHgt����M�.�?��@�G�$j�`9(<�mĪQs��@�FΈd9���������ny��Z3K� q㒶$�%��O�'�3��j�`�5�1^!~�n����˱>�㜵|����z�/gb������ŀO���[�E�:5rz 8�@�\�	���̂��q+���V8-iL���}��_0d�Zq��+8�;���jlV�JV�"��e�K|0�f��M��<&N���W��M�:��:�}O	�"}� �ߦ���k��:.�]���uo[�E�8k��q�Y<�D5���(����m�uv���������(����_.�B�U�'��+�<Z�S\�TL���c��5����}0�'\����p,p��X�:���{H�,> �}A[�(Y��钌t膜�kh�h� /�/�e���E�N�F�gj��i�a��r	���2���:�Z*���i�r��ɖ�z;���2���=��
$W��3;�:D�AQ�����B�@#]�(�n�^�����V�2ߏW�X�����Ry2M"g��X.����!z)A^7q	����l:�eW"h�z4V�#%UXŮN)w
�ȍ�M�b0;6���������H�}�f Ň��:]Xx8��p�v�5�޿*��Y��
L�>�V�3�]�Og�d�I���4�X<H�8�K�"��5����M�^~��ɿ�)�7� �>���}��4�~�li��z�DZDa� �����D��v�$ڰ����J��$
@+�,_���*FI�2�-�r��+����t �Ln�I#�EW��Ruy�y�����*�:���l`vȲy���ַ���	���($ŋ��6��ZB���w^���C�В1�1"�ts��$e��D�ں��zm#�S���x���f>�b��6p:�er@� ~�P/���p���$�	����o��G��ΰ/���P�9Kt�X|q2�gd�Y��MC�8�����y��-\S��rf��(&������/��6��EɆv+ݞ��W�I�O�v
 Ed�曐��B�� ����)[��ٙ�?�--���$;��p�%���x5��=���ؙ����-��𓮌CrdOa!�aT�@��߆E] �7��,[!�	r�e+7�����|; ߓ�0#���;���=b$�ǲ��m��+�M�͛���"i����d�|?OE�f���B{�ǳFk ����8��b�����i�l� �暓r�_X���0��{YRH1��I{B��y�mi�^F��N��%�J�s�?kզ��.	�8�)���U�Q��m�+��v/�k� �C�F��[�̡&+��W�-^U'W�g�i���8Y���n��H��swY�:N$���:3�_`�0g���S�Y��,\:�R���qo4L�T�������,Ι��6J-?ū����7?jA���l���r��ep�@#�\C!O���5�'x3 ��nC �Թ6]jd�f��=�}�Xf(�
�x� ��	�k��)�8W)�~�����~�Re�2F��Y�%J�l��Akvإ�|Ι��KSݡ˒Eٙ���K��cb�;oP�)���e�N����sq]9���+�7��#��n��QC�}���S��qM�D�Қ�i�^���_�o?U�c�}��w�������ؠm�ݼ]�b���d}�Gxj_�����V�Sn+����ԅ�;�Ę�F�!���������.y��`��r�,L�D��I=]�
����}�y�Ë19�����NBI���ݏ$�g Pբ���ied�
x������O`;��o�p�G�O$��.��+I�4ͻ���GA��{����M��	�`�uI��K�dK����6,����������	�a��B2��)�<+��s_��DJ��-�����٨U�[<�{�v�al`丘"�e$+̮�<,�~�K������G� ��R�yQy��|<�t�)9�[��u57$bQ���}o���P��O����a���H�G�sݙ�u�~M�vPyFb�{\�#8��)�:*�j�������/��tY������'� �{,�L��>'40!ۧ\�5/�y5U��3�U�݀S-��m��5M��|o+�ѨN��1l����0��I���Uc�TR��x4/*I���)T<�t�A��lWE���0���|�O���a�әs�'�2	k�@$����Ͼ�����Q��2m^y�<�h�S����$�7�ϡ��c~���� 2G0�f���KG���V��,�֍�8{���t!���sI:�9N��t�>xf�|�チCA��P��ޛ���i�В>����0�n�3�dwۃ�A����:E��,K#%11zH�[Ƭσ)�ر�!�2��}��z��pCdU�Ӝk�C���1*��wec$���?l#Ԟ�/���}P���2\���6D�NT�g:U��I���|l����J7�C|����udy����׽�<u��ML�^ڶ��=�[w�<t(�3��P�����b��1�b(__����	���N~ۦ"�������lf�؛�0�綴
�v�f�V8m���*/���d�{�T���H`�Ua�^�>������h�D����'���?-�6�y��Ǉ�<82�Yɣ��0������F�3�p\d��30S���i���֙�Ű��?��,�ބ�����
�3Q��*��9�^n�q�7 �N��mf��֏t�˄wp���~ǣ�L��#��V^�X�� 񸇿I���BbX�y>NO`^+-q��m}:mI�q���8������>��-�v���?yG��{��/�B�lo	$�a2��+b�Љ(@�Z%,�����Hj1n�di8��V�;�@�~�p��RC�}o1�>�ū��X�ҍ��ꥋ��Ai��� @�án�m���uj�]�<iz���:��X+�e��f���a�{���~��o9��݅�n� �im,�~cN���:g}�N"�S@���	&�!��E9���^�rWg�n����٢����*�6jƁ�S$���K*����/fﳤ{�ă�
OԳ�}�����>Z/S c�e�q��!����A�9�`���
�3��������^�_��eZ(pޣ%c������k�u&�}z�
#A�(ՒR6z;2�h����?kIdE�ύ��R���BC�H�\5O�~�r�_e�@���Й<דΓ����s�p��|
����I]�q%9��x �;z� ��U_���!����{�����~Q�R.��Yz��Q-=Yޘ�P*�;|��,�Ϸ�YA0�T���N��K<��
ȭ���Z,�
~4b�0�ъ&~Eý��g���a�Y�H� �
��Q��/�ed}�4bɘ)��x��m������;%��{((]0��?�@٨���UxZLt�O�+��"�ՂU�^q��!:,�}sH��B��w�#c$�["��x�d�&�UFSk�k_�?ͤ���T��'�����H xx4��8�I���ʐ�<��6/j�o#o���}��u(0�C&��q�Y��4F	�v"2�h����z�7����+��:�tvt8OOȆ��%lR=��e���2�2ݼ�	�o��"K�q�r�H:�`I2�����C��629l��9׈Fqorm^�X����;�r�IvX�i��wy�����H#G���zIZE��-����*��� y��t0�[�u��� �(E �����-v\|)�1(���t%�bN�I�џV����d/#>�����*���)<Ii���W+�I�MĞ~�U?�"ŚFr�����u|�cC.eμ�K����D	[�,�F�zM�vV�� �R����@��.戼�V"�������1�bG�o֑�39F��ݑ���{%���Q���}�V"�T��=ysq��(y~I!G�Y<���#�^�z� �TN��@۵�����������|6'I��rJ܏$h�X��g�p��|�wjC{jVvl�����#��t�k�(�dt#�Wͳ݃�t�ln����qF��!/��$�L�NtJ�ٽ@����OڣGHT�Â*���WO.�?��= 1+�4����
NAb@۶;J�;A�!�X֑A����N��Mo:�9�q>���Wy�����r�<6�gj���+P�r��=�x?'�{EvU̙���pjB�V(���XP��k��No�	!���~���p�9�^�gA��zl�3? &��^�����x�S�k�z>��#Ed���������G�_
Wo����P+�#�E�Xw�I+N�|��H�Anr�wL@�/x��BJm�e'd*yy#���d���ì.�j������X�c����[;v��Ht��'u���=�*@R�rPb����z@ֳ�)܁*A"���9�*4)��D�n �;��j�Z�K�L���9��>b��3:-�� j{K���J#^�mz>����u���͒;�Sڵ*	m"�L8T��#-�%�����2:'0a����\#�wT�?�9�����ݍ�U�uůs��$����C���:|[��j�P��釲J[��ሃ�ѭ�-8.�p��Y���n|���L �\�
�'W8�	5'I�l�o<��������At5>_QA�\�0�A&/���6�	�Cc@i��3?c��q����xR��P.�[u��f%gཎ&6Z�[Y�0V�Ĺ�Q
���V"zΧP� �$�F��6���,o�0��#>��Γ�����?�-�R�e{��-.ƥ��!��S�N�H��J�)��d�,��"��'�ؐ��}]G��,Tn���(�SsƩ~��bV���hW/� �����ձ�5%����y�W�[}�>��w��@_K�\��+��� @���Oo_�����UcE#���]��U]��d�z3���q�w��!�ЕG}ˤ1�$+}ce?��ն�ע�|_�ϝ/�e�cJ_K������"��x��1����5z��>t,��RL��-��dcj�loT��F���7��� /���g����80=ޛ��EU��?�n��F�EMӡM����^�GA0y����s�6`��(�z%�g�V��@�����3F��o*�퓴��#��	�o�����W���$�6���п��Qy9���cd���g�҅c�F����|�B�  �v������17�0�-�1# 9�Ho~ɦ��G�qw-�] o�$k%��['+S��Z8�*F��)��ށsjK���1��!�Y� ^�sȶ�#٘~�!m,��M+#E��֞�������#:�E�?c�*���~ޞ�f�;�،�|�Q<k��&���4m�rrߴ����ǟL%K,�p`@��W����0�R|��r��R�BKTg�[[���l���5( �]��v�&�\���u�Y���>�{a|˩g2�2c���3�=3���C�R�^q#�C�.�Ԛ��Ui��J��c���\�~�L-�c�C�����(� ��2�;�lQ}|쎜�*���ऽX5�u!��?�o���S��E�W�* t��I���ek�2�+��V�"?_���{���;�b�և�OK�'�Й�f���[����A��-ܞ��W:�كS<��/�^���Ŋ�o-P�����ʬk��0���%x������ڧ��AY<�
�����=NR(�@��AX��]	@�8��ՒX�M���}�M������ǉ��+%Z�>!`�U���	3F0Q�k��B�8t����C��N��4!6��ͷ|�f����`�?���b���&�F�Z0�ƀLd�L�	7�AZiÅ5�ݖ���x�
�(�)�������saEg�zMڭ� 5FW��{?e*,7�'�w�n�\nZ�G3�p�z���7��}\��R�r&����;c����g���j�Cd���S؂>�fώ�������m v��ߙ"�Yҳ�O"�}�����p���p.]N�O�ݯ1�k�7S��{�ڱǏ縎�R�Fn!*�97@I�m?�ͬG�N��g�D�w�o^B���(�ND�G�wh,H�}����R���H�6�<�D������!�|_i�s�Z��l���L]��!b��qx�F�I5Q����>x��~�fX��_�>� vϹJj�{<4�Q߀+��Enָ�$lx
�[�P����#TmbK��g�������^[m����'5��9�MsyU'����T��α <�@��ƈh(�Z}�ƿ[o�^@N$�)�vgmpff̡��1�n1\�C*�f��k{���᥌fZZǠȻ��<hAʦ�^0�R{ 鋥!�Cry�"^:��&�m��}S#ݬ>J�}�d���q�pL�����S��@q��i�X��)ƗUHKvJ��f��Ŋkb-m��������UM�мU��֦]���.��o}����ߨz�(+D������ [w���!�~h��X$�����#��@~�*�w|(X�Cw�bo�њ�wn���g�����S��t�Z�R�؈F�H1��5^��D:{b�O�x��*2�H7����f7�x���9yL	d�j�e�2�npP��%�C����U�a��c��ٕ���{'6�k@8������-vS�w��ߤ֣��	"V�����w��Q���=����R4pB��UU�2͐y�J'����#����(�l��[�D#������6�v���I��#A�ǁ����4�dPة��FIi\~�Kr��� �6��"����e���<�Gx7J,��[�'���=k�)78��m��L�yǬ����z:A2���d�8�l�*��b��91��D�J:��-KU��i�]$�W.z�;�4 r��_��)#I�A7(����.��K�[N������y]��F�!��3vmC'� +E�ձW��&)�v;�7�k)46'@\���I�g7�����
��m�H�Q�]�ȫ�077m���sjҫ�ӆ@��r%ր�R���Ͽ��K{2�~Σ�@�&8�g�P��R����Կ�.�S"�i!��ܱ�F;�k>����kM��EҘ��Te�H�Ft+	$Pg{(osS3HX�XZ��{C�|��$��ޒ3�~��G�˔���I�3tA¬���qGr���iyS�(5��,G�vD{3��f��7���o�yCږ
Bu��1�	��KUt��"G��nI��nYl�5t)�F�ɍ��p�xQ�p�7m��c����V�j�m���&:����v2g.Xf'�9�u�f������$��(A��k��[�i���T�d�b$�+<X%e�Av	.�M��x��P�Y��#�k8�3�,��Q�9J\ﯨ4��FZ�e�X[Np������b;��;�>�2�Ê�|����=x���gu�\/9z�U���1�ց�p�vJ�蘖.}���r�h0���Z���U]gO�2I�V����:jf���>��z9����~�'Oz`p���:U��jvlw�VŲ�y5��̋��'}
t-�n��ڭ��Kq�T��:	��ٓ�C v;ף��#��7�˙a�B��N�s�����p8��>y�g�ij=��Y���B�-�,�����cB�X�,f�Z����V:h �+)��8�%4��<����H+�_�J���҃�QH�y�G�rȆ��N�难j�-��]H��h�>����rR����O�'�cB�6���_*ttY�J���F��L�k�s8;�@�]��`�*�!G=�-A)��e��TG��F�cI�ｪ�R�Nэk5��p2��=қY��p`�i���퀁j��qa�(	�|õ����v\3 ���$,lgl놊��:=[�ci�t�!S4�Jfj��i�FA�_	�6D(�e��MshOs��-y��P|����:��-*�篍�Ʀ��%f4�VEy:_]�|�a ��'_��zꧾU�!]�4��`/���r���G{Ji��%�U��0� �wѡ�F>�Pp?��|d[�'2�Z�7p5��Is�7�&wp �Bq�<(�nY�RXlG�#{)Y��A0��ۀ���1j�שGS�!�&�裴8�7�ʩ��uɊd����4d�䚾
�ɣ=���
eN8����V�Rȍhixo���B�����p�T�fR�_m�iBm������E�wM����^����:׿S��U���gK�~��d�oA.��6< �߱�R��.�Mѐ�A�[0A�5瘐�~	{��49	z/��0���jUO"�[:q�g;d0�5_�in�/	ô�	,c��a�2|������Kã�>;[�Ji�y�#kAN�8�ڌ.s��:�Xѐ��HM阝��.��8cX���%�C/NE�� ��x?8�ţS;b���U$v����3
�`]��N`A�e&(ZF=�`Io` �Ί���Z�p�?���̵���-�xI�G3�[����!�T仲)�9�ayk�r�/�C��@���8[p?	jE�̴�V鎧�dI@xd��` �K��U��(�J�vM�͍j"��n����-����Fv�X���5�*�4McPō�0�8���g�ٖx%;�M+{�a>����J*'�QU�Y�N���u�� �O��rSX��(����������g�S}�>����"T� �� �?�dv��}h�.�Q��?�H��qT�3F'^fS����
�	� <�+C����@�;��B�X�g+�H3�]=���wT�gwڎ�q�+�s;�e.B.Y��a�$<5�t�-�Y"��Q=56���C�Hp��"b!��7���f���[�Z��J��W�2N��p�f�5��Wsa��rӆZؓUߵi=�ɵ5�r���%Y�s��wŁ>��_����YK�tf�;�HKlJ?ȣ�S����/s��03��/>�Я�o��J3(/jԌ����w*t�(#��{Eߓ���Z˕٢9��t�>z2��n�L��餷���ɒm��e�1tN��P�
��h�b��x�J}�u&,V�&�|�� r]���S����o�Q���]*6d��O�E#��E�*� �ST g�t�h+?$��F�G(�	�L+�Nq��[��B! �(t�c�Ŏ�i��@{8����3.9����M G7� 5-"j�0��wdb�9*紽���P��:u=j���4����fR���W�I_$|�C�{�B�E�M���D|��zH ��=*H�	O�p�Z������Z���"5����|�n�ۘ�P����x�`�Ou��oǻ�=�0Z��<V7���/H��Y�Cn���u_����8�n�]}<������0QJr��Բ��zi�:ۦ���Y����>�0�Ω��-O�H��@��"a�Ir�� 5p غrǥ�����E�`�b��ޥ�M��eM��!J����Q��K�` ��%�O��!��,F=e�r�';s0�3/2�E)FP Y�%�]�N=�(h%��F�ُK��P�8�h�Љ��r�L��q��Dx	��ON�9�4V��fs�C����㢿2(v�2��\Y���ܭ��H�W������u"�r��~�k�Z��/����$���@�X�}1�ΐ�'��hh���v��+w�+F��se����g,v-��(�t@B��iЉ������	���:��+r�֡�8��e�S���Q������Z�?�nnnW��6�)�4^��^S{V5�gj�>p�.��W�� �M�p(��b��@� *����/m`�)*6��e�pC�o5���43۾}U�<� ���g��0���U��K@x���	����-Ӿ�����Km(59A�=�o��~��a�����z�6{� }�˜���C�	ת�`q���C���-07��IJ�R�J����Q<��.;$�Y�m�4�~P��IXJ?��;�
k#79���1*S�Lu��r�Z~A�T4��'���A�)�1U�t(�������7��+oS�H�����%�B���Ϯ("r*�w�i��-�;�a�i���E|B���tb[�T+4�\�Ҭ�!���{�޿;Z\i�XyF�K*�B�Ɏ��6�Y`MU���X���������i)v���I�Cw�K=�^�=IL/5���lq�PX�\yk�Y��YP/�ق!�\�}�Ҝ����V�!
�s���ܵp�������:.Q=w�@���{|rGM�9Ok�<�T�켕Qo�~�޷a��c�M���
xH$ Q(
?o�aцH�LLg��P���ioJ�7��.8-���˹FEd<����haI��W�B7�C��@
����f��	��X �;���vת�ti�i�B�\t��LE�9�Cc���L��po()�����VK��J9s�,Ul9���\� ��V^\��T�(xop[����.	�`V՛&�a����1��d�q�y����[����I������T�s�8�|>��R��|I*`����j�u�Z��/
ΐ�^�E����ໆVX��/8KzW˳v�b� ���ҰhP�Nꪫ1b�Y�#L��j��^y'3�buzN8�����C�V:��¡���לx&ε!�TF[�����B�6G�1����_�"��V'�A����c��
�ܐ�N�$Ѳ���h T�b��@}��Թ�z>0$�#i �W(�R)@��R�G2u�k{�xC���*9��K
��z	���EJ��V�j��n�ʟ�5����	�Y�Fr�E3;h�{����;��(w�t��o3�=�8J�����j�׿�N��+V��]sc9��]UE�%�c%�SW<_����Z�3��NY'��4���E����;3��6E��"
�Ɔ�n���'^�G�� �|#&S�3���oHB�V�E�:	WJ�F�N�l
osV7)����m�y0��o÷h���ghS^�[w��2�&�C� ��m��}��W뒌�D�2&�(�벼�X�� A�6 c�� q��cm�
�4+�H͜�
I���6ؒe����v6����)����tX{��d�uu��$Z�����۬*=�F|��i:��A��8��ޛ;�TU>�k9��.F�����sP�&!ր\6i�f���!��:����=Y�M;z'�=�T=cC|��:���G�[�1j`d]֐�:y�OׅZ��H��K��Z���c-Tu�D܀k��v���%��C�E���1_;�)g������1���!Hq:C���BB��x��#�!s
^��Z`�L���n� ���M�`2w� ��}	٠J��i�b��2[j�C��2����Eb�����^Ae�5��P�#�[���Z��?��=g���5�+4P2�����=s���hx��7 	�qDe��_W぀�c�����!�&ΕB�����v���=��j`N��e(Z���k���#�nK����Ys>�^�+M�,���������$$U�x!F9�(5������m~�SE��
�i�F�� �ԞR�zj�R,������6���%!Ý���ŗܻ�������<���������=ZD�yO����0~��C��"�yƍ��ȡb��ъ��[���W�˔���Vu��-Ɗ)ҟ�G�G����65�)=B��cl����M��bh����'l�
��6�G�u���;��ٍ�1��]�-!��l�T@��Th��g��ǋ��s��3è�H�6�`T�^�u��/A�9��)h�88N8m�Z�`��WS��8���I�{M�}��><�<ӎZ5=���vv�n�g�G,�Wv\*���Ƽ�a���T��U���T�d{:c����~�A���'�BH�D�S���^��uv��A9!���+�P�"������:9���עC���*b�Ň>pخ��=�N�� �b%���F��#�Bբb��-�CN�K+�qMC�!n1��� ��Dq)�t04Eӎ�5��_��5ϡ���7)W�� �r�d�|���l��~��]v�<��h�ڙ��8'U�
9�߿��ol�
�� ~2ߵ�L�C�PL˵�6 �N^��T�=���T�&��C�|i��fÀB��\�M�06��^Y�%� ��W�T��g�CSR2
���H����<��l�Q� ���Jk���������zb�,�Ē)��W��,����d�l1i�5���s0C�5h6:b��f&�wf"��J����N���B�*�3�	<΅�Zi�����2�M8+��y�v�T��󤼸�$M�xQ�=�{z'��<L5��̓%��	��^m� �^�ݹ���5��c"2�0'�౥Ot�)�ћb�Q\BC�tm�ND�a<��O�aӕP7(Lé!�J�2x���!9>��JK\�8ݡPQ��t�4k��sӓ�Y��t���x�����|��O���5kv��}������{>x�aa�mQ��5��-�.Y���Ҏo�L�] !vO/dD^�/Jw1vKƚ�����Ejڠ�5S�c�n��rm���ejgf�;{NG���|�e�_��a�����	E�	�7�n�~�؝��D�8�E9�A�Ih+�u��aY}���
� �4��qВN]��V��T��	�@%`��|v��. ~C[�2���4�������ɪ��x�j7��knE��[m��u���0���D4|*GpJ�����7D�|�4�ھ�@�l�UW�	����6�}�qwu��?'�.�0G
2��� Ɲ5'hno�x�
�� �]�/j���E�0%"Qh_�GA�zr@���Mw?���'��Y�hB��O�!=�t�#��.	;�
��?���+����ٌ�	�l�F��[D*��l2}O�\�!��x�Bik=V� �Ž���=����{qֱ$r�(n�/�ڱK)!�B\O�bwZ�qA��~3 &`�Tꥵ��Z*4١Ŝ��i�����-V�[@�">$|�v3N:'-�y2�:	=07q1�k�_h�V�6`V���B+X�(Yx���%���%k��G9��{�E��Jg��$�80�X֡��&@�m���U�H>ɜ!0�a��_�9;5�.��"�a]8i�����g%�m^J,G8,���U~�~؝.����>|;�)��q�Q�i�=g2��U+�E���Q�:Ae�rJe_QG�	,`��C1wD��T�+SvΡ�֖�������m����r����F��
��X�2��3۝��Ns���1+�	p�9�~�����ByP���掚�)tk�z�z�%Q�k*�	�ה/��c�����2�����~�\CB�OR��&�)}R>��P�Y܆W��e��Y��E�9;���@�F�?��[�������R0O�
Y��bP����f�	�,�h���2H�&���^8GڄRTL^߅�S+�4�E��0�\�Ϟy�>S�5Z5�.q����$&e�l2�;���t�QM���t�v] �Hd7}�\J���x�!|�;J��f�I��w�2|o5ƶ�k2P��w�^_��R�j�uUWؘ��.v��a�A�k�]�Vm�� $*�ztzFo���)���d|2�	u]�S�{���54P�͞�����J�U�}�fD��k0�������-�P�5/o�9��0P6N��s�sQRT���2�AZ1=6�.����q����+
�(no�֦^+�$Ji��?�u3k"7�h,7�OUiw���Z�Ո�D!D1�� ��������y���v���CJ�|~9=���-[T��C�j��`�β�W3Ŵ��D��CF��{8;b�5B�?��k�J��p��B���D{�~�.�;p�b���ޓ(R�z��2�CHYuC�C��#Z���i�����Ed��l�b�M:�C�%꿛{iT�h���j{��jK�T���4:^lKႶco��$�~��Ua�q��A��p���5EZ��Hm��36�ۧ�~ m��7ȏ��������iK%�&�tG@��!��ze	C�M�؄�� ׺��e2q;,�d�����ۥ�	�wl�?^N��[}b9�Bkմz�I�9_��������؊ڕ�LDV�18/	�
f��h4]4��wW�Zx��$��%��M	���ј���A��!2��W�c�K:t3<��w�n��I>t���ς�:'��ǋ!�PZ��:����<a�����".��D��NXJj �fF�)��\c�nn����w�ڭL��>�*mVF�r�>'x����5�"�v���e�­�`�+�����.eĭbPS?��r��9�n&���3lm���#"W�T�[�1��!�Jpm�DJ�Q7���|xy\�8��b�\p.�O�6�.mL4���M�T���7�g?i���KGڳ�ʲ��:xp��)���F�oF�p�b,+�Xԩ*z�@o]�ɁA� �KL;g �Io�Y�T�;����B0�$�ʯ�*>�ڋ�S��2�?t��
z�c$+�����b�}.9��[�ݸ�ގs��?%_���G=%��Y~�akK�s�����b�u�L�G6p2�r1���àl^�; ����%��?P�*��`4���L�_�Z�/�-�R�XgQ`5�l����\���
]<���)�����c�w���գ@~:�}(Ӵ�WďM��N�t���[cGU#v�X���N��pM��9o�|j���x"���>i��	]�	�s[�o�Tfي��h�� Jk��ر�`�q1����qľESU�x�k���_�zM� nI���,�����(�4���aT\����x=�'B���HF����g��!`��R��y�[���B{���q0˪��oUFr~
��q�d��+I�#ʏ���6�63R~T03⵬�䂯\���G�]���Qv�-E�	���-�����{(lLPM����n�ȵY��7>��!�]j��<9�S6���D6�Ry�M�/��W��F����kN�JKc��nc�%:m=�i�(��Ly1@�9՛^\�����K������)���2��QZ�;F:�Q��=g��H�q�72��.���Kx����K��\��C�Ր�7�w� 	���*��U�8 Y�[�:1g�iAz���V��-c�J#�/@�w�)/�� �����BQ��(/6`��!�F�:��p3ǤaC�P�h�t����B�<&�O[a��n]�S,AÏ��Ez|�����6����\�%������"/N<�f0 $~a�,�k�V_��ml8�L��SL��]�� ;&�:T��6�#Ť�P�'�o4{48��
ї�C>N�@V�B��f$G��*�Z(�"���W�c�:y:��r#���['fy)�u���� ��������#�Q?�u![ϵXM`�*��?�A��N�빛�Z�zm��m'"�샸��P���Wէ�����{�J�t	����A���3����`VZȣ�"V�����aܝ�a���n���$��i��ަt��9��ָ.��W�
�B`�d���gV���$�A0%��4�v�������ݔv2%���9*d����Ε
m�4Q,}����V�2�\�+ıo)�0����b>���N�~�[����_7j��,1���0���V��~��$ `���C+#(�=`m"��Av��k2��r:���7���:~B-Bf�#��K:y��'�"�t�`�q�;����W��wu����S�ޥEdhq,`��r�ķǨ�q��m g~*RU�#U	/�8�@�������[u&�+�Q �=P��'1�����vjM���_bO�o�w�߲YmA�SXo���)�'�؆�h������k��BȺ�j����'7e��x���A�1Pz�g�u��wS���M]��M��?��&�V�h]�+Y����z�O�������ЍPy���%��Q�?�æs@Fi0<`؟���?}��Zs�Z��0V�L�MéB�o�)��Z}߾�1s��;<Y��p$�盆�� ����K�)s����~E�}�w���r?�bW��i՜�z�	{L
��ؽ�%+.�������OK��#�N�5�����=u?x8�2�%p��RB�����(�����Z�)683r�ĝ_�]��fQ��A�.�׆��9�ɶ�9�x�Cr<����*����ޥ����F�=� ����)�Q;�]����L�v|�X��ۼis��|#s�I>�v��oH��'��&�O�~������B�nx�wX�����E������8%n��/�(�"��E�&-ek9b�E&�s���E�p�Ce��c$�����]��%F�s	�ȵC��an�;��f+�����%gp���b�6�IAr�Ώr��w�z�J�f���L���3,k�jk*5��z���WC��'�ϯ�s�6�Q�L=%����@�l�w��
L{�v��<[:u��]@�*���|��v4�5���Ά)מ6�Z��h)&�� �w{�-�ȝ��Q��Z\���s�7n�u�ɻ����XVE����Ϥ��{��l|�U��:iF�`a�>���A�k>��5��Y��$��[���<t�(�T������R{��`.
t et8��_)�6�`�Pċb�����uN�*ǖU�{�����W��;������Fg��J��a�Z8��/��~Q�$R���୬���쪩��\%eq����l�h��I�-�*ȍ����o���{������`�x���%��S�FO��@����9�@�l�Y���`X�g��l������u����-+N��d u5����q>L�C�O+Q$؋���ڣ�{�Hlݢ���%���M�ި95Q���O�����P��SG5��vϘ��c�3_"D��A�jf�Zɟ/�(fӚ��n#�C�[Ϫ��h�)H��z���*���)���p�r!=L�J���V�����#)!� K=��Q4����>R�=^g[Ƒo]������E2�`��`���_R~Zf��}Z���9*��ý�|���#�	_v�E.���?��j��QL#���.:�������,)������yf��vx� �e�S������*Ͻr�{}?ոϰNO,���s�*�D5�6����ϒ��C�A�U��46$��S�^8t�6T'7�ˍ�C1P�#�R�H�3��
����gݾ��OX���F�x�%��f3�l�$3��$P�z# ͍^�z��A�}w?����v���}
�حMY��󨨏c�M���OY��'�8]#�yU0fb]����}r�`nP=�y8�`:C5��A/D��Z��ՠ�U�,���(9����.�L3��|CI��Ⱦ�L��܄杍�rVSu@0���sxZ-%�	����`M��+O���,�{������.^�)���Y ����p�c"PY�å$k|d���ِ7'.෈����ERq��VfØg���]�R^����
DL����}\��.Î{d�r~Y3k��x�O�����J��7Y�]�q�q�ʇAV9�r�ѻj�o9�z�x׽ i��D�9j���\���`��/�k��K�/s����;	�$`�e��9APa�/m]4�mv1�*G�o�ŗ2�Mo��c�	qS��zQ����˻]T�;�Hyw��T��O��YCI�zi�ū��H���H���[�~���� ,�ԗ�1Z�*z]��Ϟ͝�*>Ң��Aj��xM?h�ێ	��-�6
�T)�}m��9�����h��u&y�<A� �0����.��! ��m��dc�����Ys��G�O��� �>���FU-�8.��V�^�Z �]�)qu�-�l�����Z?AT�[Jgc\$�F�캲'$&�jwVPGHR;�K`���PZ�~F:WǺ�Ğ�����c�~��~/� ]�����}�|�]�v~F�'���x���(;��3�d���]C#����2�z��ӱå��<�_�h�p�V~&:|�|Z�.�;N��AS(�;�E���n�D��.�b�Z�e��*��Ο�Ok�����vR�g;R��g����q����ω�zK����dE|ԥ�c���0��`Ԕι�h���,t�K���XԾݏ�f_��0)[lH��`Y�
�����k�=>�b���8�x����1᥄��E��(¤R�QrE��(T	���[b�YZ.J^��x��`"ILr{z�ٗ�ˌ�$�n�_<M��a�����ٽ�Z�bc��'NtV�s�;?Qf�����B�Ygs|�9���5�+�iu?��C>i*�p��N�o�&kB�������I�BW[ ���eRoC�cз|��;� K�>_ݢM�2Yw� �y��
}7���Q�X�Y�D�Ǆ�r�i�sP���#���	n����ȔI:Fn
��������%����C��m�'�ส��c���!+n�<��^1�(���3���kYp�� ������h�.�����&Ǳ˦�3K `v]l��0P+iE��#^4dT��&�Vi�@�y�MnoK��2���,"�Y-a��v�؈L��K����\�[7y�����tU�| Xc��(�P��8���S�{��a�Ȁ������xw��k+PSc1%ݝH �����n�/m5x��W�Kbܜ{��$������0�L�p��ۆ�4��~؂� �������?U��U/��'��||������4�8��������ZŎ�/��f��^'=��	i��χ��ƚ�IG�V14E9�ɛ��5P�k���<
ן�܍c��@�:B=�({�?��f�������8٨��5B�<u��w�o�*&�)o�J�?e�%��ړ!:��0�L��P��SF�ZsQ�js9��-��Bh�i�3�%`���ͶTd@���3M�2���qj�~r�
=��Hv�U����m�{�.�喗�#wr�	�l&�u4�}���O3�~��
D,���5��dB�{eҪ{�]��ڊY.��ʜ������Z���6�-�� i��7�.C\���h��%���?]�.m�:S�
�>\Q�����y��a��8)���4�8�m�}� )q�V#{4[8�L�z��m��.�k�����Js>f8�����w��:���Ы%KI������-e2;���8���՜�Ӆ"��U�r��B)��ӳ�悒y�����NՇ��>អh�3f�{�<���L�k�*v78��!m޳1�0կ&��;�W(e�~I�S����Mz�ڿ���F�d�;�1�l�|�w��!���[����1�%S���&��T��ͲG�C��Q?�ꮚ�_�ׂj���T$��l'��)T;5��t��c����4 ~���ƕ�p��<k�j�X�@'�i&(�5>��^���@�2�%/A���@y��"�
�_��0���<�'��i���+�(9ЅR|����p݌�r#��H�֕n� V�hI��7~ �D����G�+�a�QD��x��S�`���S����tgzc>bf�[��#����D%�C6:��=���8�gܐ��x�<�)H�,�μ����x�ļ���Alt�҇�Ī��T�<|`�-���j+�G	;���i�o�&~5���أ@y>O��s!z��Xǔ�f�&<E�3����Rv=:H��A D#I���S@��ߗDI�+੹A��}�P��H�	�>�װ� �j<1�k�2{XN�y����s�W@�H��A��x;,��y=o\(J�w>�������g�n��*�
kalˌ�!
ˣ�]q�Ф �|A6�Q�=�=4�dTD
�+��;�w���8ۆ�x�3�ɗ�5�[� }�{+�'+����հ=|~�����`u�G�"c�GK��RiM�Q=K;=x v���kh��V��:�Р������%v����c���X�xasV���8K�Y�6s*}�#D]�D��u��:��g4/?5���5��`,`�EV���x�;;{=?-�(�F��Lyv�VY��J!J�d�/B�]k?�%1�/l�b��.G��q��t;!���t�"�q٤dh�	+N.��AC�w\�'�]$�i4��[�3�5���ͭE�<�f���u�=���9WD����c�.�WA-o-��k�;��ۦVk����x�tC����I����nLl��a�O���y���5�/b:�Ή�X6���<!K����JwԆ0Z�u��n*�����?D���Ӆp�(��e��Z�]jy�,+ q���|Q���A��_XS���϶qV�Ky=g]��8}$�1���s&�b� �fv/t[X=	�w�aB�$?�;������[��{���;Wh�Y�gS�P�F�f,�q<�芌��BX@y X��C6�ԛ�go�B�a�}G��r�H���z{tJvM�����bj�JR?UQb@��r�fsNB�єl��|ǳ��"�#�>3�*n����GN�R��I;^r�����Z�6��Gǵ��P8p��6��b�"��%]��O៤��G"IRR.9�;3kK���s1��t�/Q�߼#�ѷ��.	����v��k�?C�`��D��Иʍ��`M���I���m��Ѥ�w�Q5�JYol�Vd5��[MuVb�[[���J�:���9@xkY�(�S�F�᡾Z�=�EU���[�gɬ�R%�p�c��J��l't��?A��~wΤvs�H�~�^~��D����G=Fj�?]��6�巧��J��:cYgL�Dow&@� Nt���a�p-(�(�x��T����n��������&*Ͱ|��`�V�Ԙ#9h����p�N�Uٱ��E��ǝJH�^�a���?�����߉��Dm�2!6���r�����Qc(ᯑ	��^�>gQS�|�\�����,Md�����j@�|��8�f��s&���򑼲���:��V���W@mB�O����6H^>�`w#�n���&�>5������~������s�6M[��OL�n��@c��^k�r� v���p���7-չ����}� $G�?�2�A����C�ʈ�ȕw���/��g��l�o^�_��1�@}����V����e�B�e �"h�#6F�Q{�'�=y�����R��B	�EGC��2�%(�Y��跆�DGsn��WC�o(+��\�@��z�:)��{ �������=��:����ә�|��ޙX�(�I/,�wm�X�DBq���>M�Z�D�"v�y�K.�RU3�Ƙ#;�f����O�*��%�n�Hb�R���(�_�
Y�&�B�5h�w���!�����6NX?#o�}CK��5�f�k"S[�z���ˋ�|�Ϝ�4>�i�,{�13��nHO������Ik��n�'A�'.xo0�1�zB��3 3_��E��mG6�	�x�4����x��^�F:����~%<�c"��(r��b$4�����X��u�.�|+�l�[Ej�K�t���UO���	B^�[aЅ��ކ_R�6\�Bgη�m@x��|h�gٛ�}g�>�W#ڤ?U�����g����t�ӱ �W@���f�nD�a��96��,�zΌ�eK��|G�@W/OI�S��"$�Uobj�g31 ��fB�'ٮ�K+\�8@7�T���ov���j��z� xT�c��_��F�8j�N��hT��$�y��F��ϙ��G�S��Ɲ�i��]y�/ �"x]�A%�17���PNWՖD�3�x���0�I��o�<�e�C�Q�"%�QE����E5��8�V��u��ڢ� �2�	oŌ���=��z�Υݐ3�q����6s�b� *�����S���?��F����SZ�}�離ȩ�[�:�����Dv�'fna�wĐ[ ,�#�R�]��"��
�m��,�*��B��E5V�uT�f%��u��wwgͦɒh�|�;["ɠ��Y���|�3�1Jc�{�[}���1��>�(��Z��pBX�G���G'5�s�[1��f���T���+�m��F��r��G��C��ä��P�Hׅ0��`������WJ�ulu֗���������I��%ZH�Q&-����©�\�2� M�k	6��n��r���Ք�O)����F(�%�A9t��sV��A�����o��/le���_���ڦgGڐ^H>����+ܜ�5B����|�ʢ�f�wFD)�9�Ju�+	� �b�%��;��>�g��� B�V�Bw+cK��!��Vvy��1�J��������Tm/�Γ�aԁK,�D��1p�����2Ѝ�}H���C��
�tnM�f]f�]r�o��^��.�A�P����boa8q�����L��\E?�K�,��R�6�E����>��y��|�6#��"��K�a��5
`c��̼,ZFYfzh)�N���XZ{���[�Sl]�"M�j�Iʑ��9�n�N֔�{����K]��q�4�c⒆��a�^'+�E���{RH��QW�r�(�}�oC���:�%���=@_/��`�g�����s�����	�����Ba�"�Wy$�Xso<��;���a��ϔ�r�Rh�&�ڜ��L�MV~����v݋ �����g�8����O]:\����߸u��&H�t�����Iz�j�{NB�a4x-N��*�T��mfgL˨*�fg��QA�%��0���oq�<�sü:ڍ`� Y����U�9�(y�!B�\F�B���@� xU�|򚋙r9��>� �+b��Wv[����v�����$,M��I(?~3�㷐����ӣ\�퍽(���Ha�]lO5c�FcT��>xp��@ �dŤ�\3t|�,u;�~E��7Լlk�B&��٢���N2�#�g�D�/�9�@�����d{ύn�O/T�-Y�Q��j���0z5���b�-;2aKW��,�,,��F�������@�M�T"B���(/�?&�� 6����_J3�ω��N�Y��o�fM�;�^�H��{�W�J�?�Q���p�����n�2JtQe}$r_L��±��"�� G�0	��K+FIcz��dƜ�CbM"ם���	w9����B���k�Lʷ�T>x��^ɝ����u��։�2��-ӷ���pE �������i���j����Z6����D�Zp��%*^�����L�i��y�g�&���/N�K\���T�#-�=�h@��ɖ���g��&E�Qɳ���YRe���{+�̏�n����Ȓ��]U0e3��,�^v@�_��=�sd�s��R��x��H=s����,��)�7TQlܯ&g���ӡg���и`���0��6I<UE�$�K�ӽ�9 u����KW6u*\(P��M�����Rg�0�u4EFHU����H����]�c�U?^�zf(X:�MA����Ξ�	/��
o�%�3Dn{P�֩��jD�O�K�Ӕ0�?p��3��rSeYĿ��D 6:��л�b;nU��}GL�I�7S������C%A����n&����� w*C�h9.�"]�U0`�f4����~I���F�|���}�	�r�r��t�w�
��[׵u����Í;c������V-өL#\]C�߂q��r=�.j����po`�C��� �U;� ��Jv��fP����Z��
aS[�
�1jۓ�Y��L��e�M��FBp.�?7�z�$[��Ź�u�v(�{��(d'���;Dw�!/��0��O6�RL3S�B�_zZo�5��sAN�����B� �[�G<L�ʪTpHq����~Ǧm�7��-��ٽ�0*r!�C��ZV������=�����B0����s�iEΊ����y����kψG�@K�>�Vfߧ�1ԭP!z2����d��zI�T�OE�c���H�~���qq�k���<Џ�@<Q�4Z&ڳ�����,�:�ˢU��B�Ծ�\<��=$���(."m��x�1��0��u�Z��yW|���el�?�#����u�Y�����7S��N����m_ҝo��vڷ-A���|��e�CLs��Re,47��6��]}��ϏzI��Y3Y��脍�����]'�GMG���y)���k���!nNhE�kVְׇ��o�*BD8z�>�K}\'3�:ڈ�k�:�#��P�^kspRp�bd����t��*仛D�<\�CD����ާ��{��l���,B���62K�w�����AU!=�}��ҙ�2r ��˟g=���F㙜���7����w{��f�]Ҫ�057dx#�"�rt�̌��$k'��L_�b�#��\5���l����I'��:AM�+tf�C�Qi��iK�����Ɠ�i�^����o�7��@�pz�\��rs?>�qvֱ0�s���zsp���Y
|ekS7��� |�ǜ�/�8�ͳ�P}aʟ�ۼ��сG&T?����e�
J�̈́%�,\o����^U���i�?�:<�,z�غ/�N �L���yΦ�͘2NȌ�0]1#N���+*���*�m�%=��t� j���6�K�������I�:Rp�j,W_m�7���;_�XZl0}O'��y�|�p�1v|�$Ĉ�:��	�z���Q�������)�h�1��V�<�f�G>�O��"7�׆�8���Vc���0Ļ��I�:zÌ�(C��瀲�J���9v�vb��&Dy|�Y��ݣ���`Wu����~��R4_�K���8O����$�,7ď�o��I���w
c&D��]K���b��.�Bv���Q�^e</CBB��#H;�18��Q�K��/�w$e�L��L���1ŊoE�F/g��|PS��ၙ��wc��7I���3o@ ��	�J�A��1e7d{���N213�!�]E ��B�iY�Y}��>��,���	��s	���o��(���
Ȼq�5�?๞�4j�A�+�:�G����"���v�FMKN�Ӱ	�v�t+�H���Z/e����F�d�M"w�9�y�@Bp!/�Ovx{��#�Z̓U1��+4�V�^���=��Uw@���ީE��\���
���[s�Q��<��3�2Lz{
�F�%fI�����;K�u�`=�J)8�6�]�����6G�s�L3��8��mr��<�ux�ي�mƘ�$�k>�b�]��+iX�*0���_Zr���_��]#ԝk1BV�J����p�W���zo�O�cz�x�QE�S�@�_=i:I�؎�$B�pg�zv�[�[�쩛C���CY��6�,7�=�J�"�[/k*!��G�W���_�4��*���r��M�'ݽ�%»D`N�ͣ��	C�y{3�4�V;�ue-3"��9�+��B��H��l���Sz�����u�N�8�l�IZ1Ⱥct)�$Wo��nlm �
�%*_]�j�#�T�vr�5~��֐������>�6����z��"��%%����s���&Z|���~�U9h��I(���3�`�'U�h�o���)�z��' �Z�8ExUg��c%bjz���sr�����:�8w]3�,
��]&A�EЅ�ا�)��oU��ޜW���[�tXϜwUAk�>�^2�%9�\��p5o$��r{�e�_��:�!��d%',��P�^�v��]���a+p��_�ڣ�ߞs�>"ig����7~K��_���ޠ���3�6};�#}(�}�"Ѐ��DgvWR*k�'Xj�@)�0������S���9��ι��M��M�})e��Ө\Ӗ*�)E"&��r�n���;���[��/?�3Zϙ�K���٩��!~G����e�%5���n��iL׵��{5R]��HH�e��$Q�:��&�<\���ִ�7*t%R������o`\�ב�e[����0��d�O(;is����kx
��UTZ�mb]+��?�D�|�L��!
Ӣ<	�g���V�Â���c�/аx�?o���9�4�>	��Њg�5̆��g�A��Q��MF>�KN�M�Ƚ����X���z�N�ʧ���*�΀W���!����d��\��򡐸��l������:y�>t�	��e�%1K~�o��xYD(#�Wi������nHS��0����t%C!���9�@���V�/f��Ƙ��Jf�1���š�	nޮ�����#�I}�� ?g����X���/Y"�pj��b.��0�նR�Ϸy�Q�M��`uZ8/<��a��E��9T9�����Co�2J�q�� �vL1���=�=۝&/&g"��	���&>�Ǽ�R��ػ4�4_�q�~�q>�#*��8�4�S'�-qX��4��~à�4L�|�<=>U~�����ӳ���9��G3𞂤���鋓��~����z�R�����=��n��d�Gԗ��]>�!���D�xn���\��)�I�El&y�y�]�hAi'��"�T��"�J�[�Qz��x�U�5D�������k�燩I��[�hX�kYQ��R`��!3X�o�qI8K�N�����="��av;'�t
v�c8��En��Ba�C���;�b�T7������^�+k��s�ut<QA�����	g�_��%�{��'$7V���W���v����[;�:`<z�A?����S��4�����(�A*��o�1!΂�y�ɯ���W����&�m�D�G��"�Ƀ���H%�07۹���e�Q,/c�����P���@|�+;ͯ9��=F�I5=�a!�׶����� ����$�oV���P���JtB!�%��- �F�H�`�?���=�����T��<�&��x^o��THpO�Sǫ:�	�->:�.� �����&p�]�7=����1���i"|������$[��c|Z�#�f������YY�����}����PP�s�Z	��j>��`�k�o���k���L:�H�%�~ܫ�F�ȡX:)u+.p���I)Z~؈<��UǦkP�ndh�I���B/���r�ꎮ��� )�^V�p8��Y���|-'Y(R��3�u�S{���砒����y�:WtU��ub�^؊&a���!�=$�������`o��V^�����3������*}Μ����e#�|c#���gHLo���Ij�|���(�zͶ�-r����7mU��	6��Zr��;���>+gĶ�Io�����.�9;8�;���Ѧ%T���]�&	�Ķb���ʬP�����@V��[��E��MF�oyD�*��i�u�@�L8�
cq� D�;��������?/a��?\Z�G�(9	H�H-4��$�^��?���ì���'��3�Ȯ�4�E�o(C�ul$�Z����'�g$��4���s�*���[8�/q�D;�Q8�b�3Cc�̀�7����d2��O��ܐ&L7L��G1����8���iN��e׺�&�팶��`	L�,�r^>Q�Fh�9Tx��T��d���=G�s�~������@ڄ��4�D[K�]"��;��������ډ@d""���t�3����^���ϥ���Ǳ��{�0rgfF:�gA���}Dϸ�����{Xj'�5xR1�����Ix��AÕ|��$��L�����'{Rc�?AB+�2�l��ڝ�3��*�ĵ�g�����W�1̢��m�����f����d_��<.Ӽ�ڑ�!��Ӎ�z�t� !�f#��zp����x��� X��cr����7C]�]-���F�$7a|Yc��ԭo�A�g��'|�8����o`���b��=ye�� ��^��y�Nun�x�z�C�%ʙӺ����Rz��̡K����|/����Tj�m`�1W�6d(��k�9�H��ђ<d��"e��l(W���w_L�ۍ��R
��Ҕ�nw�JX�Y���0E�pj�������l/�?��K��0��2')��(#�	(���
�n�k:!�{�!8��%Y�[ߣ��=uDý}6%�K[c`߸�
h�o������Р���\�z��A�<��A:u-o�����\(x����7�pA|8 �(�	M%�!��z�zđ�3�k�c�<�[)�(I�8�G����*�y�	Ij�RpG]/��>�>��8�(�ȅ��A�3ʎ�4�4%~�Oݥ���{���I����|�X�~��y�q��H���9��kV���
���m�Ơz��Y��P�H
��\��v�%{�t@�VVG����"���@���y��{e(�M2�1�X�>��aHX�uڽ�8��Ѷ����T��w[�M�dU�7�U�1�v����jjNn��7��4��W�a��N�����X�k2:\�K#��?b�45���	�u4bC�N��a�	���ȹ.���,�3����lO*��~�%̮QIg��/gZY*w�BE|,<G��Z��'��jC����,yp���z啐��qg6�� U^6�#�|aE�K��������$�>?����v�QF�gG�j��>u��?�sjY$O
x�?i$����\{w=F�<�$����_ieQ2�BΤf���`w����	78�*��^Z?tM!H�N����ˆ!��%a����ǖ����༠Z��#6������7�����"�(́+�s�f�������fX#���{r���o(U�ۊ��iCo`��lę��*�#T_�T���F�2v�-���1����ω�N[����p7?w��n4u-���f��\Iy�4�f��C҉�Q�2mkPEJ��Q�Y�S	�����tW��Ge֏����%���œ
[��h��Fr�qZA͝�8H����EP'N���U.C� ���������Ch�|�H�Cթ�h%=�<�
�>l���i�����
�.��R��̋��#Bu|*[�`�/����Y�<�6���z�:ٗҳ"��Vc�q�6��+�3=ܷ�y�0zs���J�IWl��Q���M���c0����X����M�9�$�77��&���F�X��89��a�l���r;k�y�/�|�$���g�o<y8{VLI��\��K���_�j�~=�e���f�d�G�傘�����b}�(�糭B1��#�BL�ly\�KqCMOt��u38��
Q��o� �8���4v�<����瓝��Z���p�*�����=b�E�	��x9��]�(����=pV3aMg#��=�E��l�}'�-���sf׭vlp�m(�3��e���8�6����j�h�Kn���q�ɔ|"َ�+��b��Ѵi���1N��yq�˽U	$���c��.����o,���Þi#�x�NO�c���{��e��N��ٍ�W0>':_�um��_0J�ZCo�h�A������(	��`g����{�rNZ��4�+3ֽ�U�?[�;`	I$��m�)R��4j�$��՚�֙��#��I>h�O_vv!��"�E���h��k�D���7�"W��)��>��7��u�<B��%,�r����9��/���e�\e�����Y��D9D�"-]��/{��|�MO:]�t���4R���Y�q��wǎ�~lf�j��ҟ�d�n^=Iϖ5��4��
�w��zr���G�8,ݝ��;�\E�d*0��zT(��&����ZS��Er����{C��Вn!zFᘻ(����9�ܽ��Z�,)�xz���=��P)�m�]�nv�G�c+���R��0�0%a7L�I�O����x;oU烲+���-�����c���FCۥ���;I��1��T�WG���������8B� �4E����V�.�`Z����8t�0�����\�W�1���W�+pIL6���5�Q�a��Vg�6��O�K�)ms;�r2�8�[r�&}��g����}��H��=��
��h�����jt��(��cO��q��W6G��M�O��f\�+�js����*�nnl�ҙ�i�9��e��x��,���z)75�����f\�KQ.P��ѶʍX'?6�E 0 ^�f=ِ�c��S�`Hܐ.ZE��x��S���'ߔ�%�D�_�B���Y�нQ� � 
k�l��&��B����K��5�;�euO%X)�g�'nsCc1N��{s��%hs�^�5�t�e�a�w3�n�%�+u+g��}C�}�/oԛ����8y�z f�����U���P}zݻ�Cm�K3�r��O�:��H�:Ə��ǝM� |���O��vFR��v���
�9�)逶��T��8E���M�2a6�b�Do��ՂސPӮ`��Cn� |;��J$h^͜ǽ�8t�ښ��nn ?���6{���֦�*�eg*Bx�5lt,:���'sw)�5�E<��B՚մ�>�Y�1�$�D�+sB0��D��Ǟ�?;YLW�*��?�Q�a�`�N���u���(���*e?2kx��#����Lu��}l���á^Go���~�H_�WàTs�V�<�y]�9Δ��M�VB1���[Tf7]���;=P?���i�%rG6LF�v�V55���G�'��=h�&��b�́��޷����X֘-P���oA�`*�ќ���Ȯ�iT(u0��<��(���{f��2��j�h��FگP���v�i���2���Ϫ�T�`x�.�gjNV.��8��=W#>p����\���D_�g��.�{��T]坧6�{f�S�[�G�dҮJK��N$��;�M�u7�Q�NK2e�>Zq��ɜ���XO������4��3�D 2+l`!�5R�S��,�F���14����à�n�WֽE�1]�_�Pe?��am�\�>����z=�}�U����U ���@�mtC�;	�� �FPC��n��S�A{�<�2��z~6�xZ�zy}��ʷ~R-����̈'0	Ȱh/7:T�m_�����7�k|�y���R�g#��A���-�<"��(�Fe?��E�����ET��+rV�&�����
�4dU�̔�>
��`�ě�1`��h�؞��'�9D�1fU��ݵꊖ�Y���e�	����j7�,��+�cm�r�7���~�0�O���5w�~���ƏE�E��.*�l�.$����������o�Y�� 6>yp��	�����`��)�%*�z�v�tb8C�Oh`>qؠ��{��m�pS�	y�!zqe\uڒ�L"��e��������=�9=�����#�;���V4~Hx�#> 6Tx�Gl�N��;{���3��F�H�����SCfnۺq��Ώٞ��E�ڑ� X�&�E�ȱ��߼r1EID3�+a�?B�X>.`u4w>�P�,K�X�@!�f4O\&d�[a��v��kׯ��'����&�7��t�#�N�����#�M��b�0���X
�K� �w|C���:�Mf/�Έ��b1m�"�M�l��~��K�hJEt�3b.�kX�Pӥ���ː�;\��)mB����4)����g7jd(�D���c���d��7ֵ��멇z5��9�/bX�sX�0ϑ�+�}�|�^'16�Q�J�=irC�1���-+��@!i�?P�{�L�U��Ӫ� 鐅�9�b힜��8�崸H�~6��8W�j(�J`l~�ܡz~c�'�;�.�qԨ�M�5OIO�&�t�u�d�!ŔO|W&Ɨ-�N�Z+*�����v1�(׹�
�X� e�ϙ�Y'D�M�f��@b�c�`/�2J%��3t�苨�I<�Cs҉��$�3�FGf�#"������� ƒU�̣|��Ġ����b�t����KE�����j�]6�DؤC�C��_��H�_'�fH��.��P�!��-�v������9QH	��4ޗEg��OS�>.��Vtx	y,�7�&'<�
j�0�z]�v�lL4���&��2����eM�?�r�W��d���Ň:�&Df
�f�/���V6��s��&��[�C�5Y �����������p��V%(�r5���@�8:kc�����[�����5R�G�2�b� �������EJ��#��w�[�^��[���l�����O��i��:�649�*d��COT�������rʎd#;�3��hL@�x#?�۷Ww���,��f�t������� F\�Q����!N|9��l����B$����ݲ��e�c΢rBx:�R�L"�r�3�%ބ@���0�j�[��h+�-G�ʤ�z�Io� �"��q����Ȧ����H!v��V��Y�������:apc��-TXPl|o4��j4�A8�>$\��d�27m�Y_�PX���6��z������.�QF?{���nsj��X��j%p�z�H��wC��|%�J�w�9�7u�k@n�%6v��|�q���'=����>.�^s�B�]�O��ͪL�� ���^�=��'�S��8��@I�+n�ca &�Vz	뻔wu�`�f��MX���B���'W�	-	�HHh!<���u~�4���Q��{��,&R��`|�"�;==�+���:x/ǣveN$Ss�0&��_C4^�M�vi"���U<ט��������5"�L�p��U� 8@k�{v�jqP������y�&��l\��_~QnQ�CIg����Y��9;���E\z�l��vd�8�2x��-ś�xӌƧѝ�yQ9�g�7�l���W<�桗������|# �n9S��b�g�B=���1�5c��e�?�j٥d�i=u�?�+
	cU�̍�,{�(hw�+��_��Ze�l����Яf��c���)������4�`�®�߾:�a��L��&棋��ͮ�c]���A����*�JJNR�~����d��9��3)>�Vo���\B"˄�Q�[v�n��
�gg�5	qx#S�A��i-���ޤݭ�#�L��ܜ��= �� ��J��1�C.���*�L�P\�N{y���w���w|�Zqk�>�vcY�s��"��c��ßXN��U�A��U�JS��k��4�1f�[�~�p�@�'��"N$�k��E��X�P��n���M����❢�`sܭO�bux����xI�acCִw-����[S��<sͰ�?1��.V�����Q%ۛ�o�Z{צ�U��Q��r��&����'N�`}-ֱ�y�S�j�śs((ND�̸���9�Y^��2IˬU���9h���zd�ڍf�'�9P�N�f&4a+(��QA�,�1�3�P����bEq���ǿ�i�˼C� ϒ$$�ĂZ����`S7�}���>���b`�3m@"���iH)S)�5����MZ��@�����Z�D�?�)�	��$z1�f
b�V��U�AA���w��+߈F) �}��(_��e���X�� "��-dҼJ�w����Ǆ���edowbc�h�C���Tꋨ�B�zH�%�����d����1�����Q�}��z��,��Y`�3'ێT�H֙s��
s5y�lPTOk�2�5	�VXZ���A�ux��(�jry��f�+4G�'@kL�*��/o��+0?* �h���!U�:�L��C�?\.l֡it���%��s��9�H��J�ޓ��Hԇ�6�Z�A�]��J�c�Çr��a���M:/���}��mC��"�݅S/M�,&c� ��~�j�����_�rR�(��,�����$��IޙL�D�6Y��s���_3���K.ͨ��6EkZpj���L	eR��{��!��miݺ6������*|�:�QͰ�h򎷪y(�:���>]bV���߼0�~'�7d����!�9���YЇu�W���k���]C��#V�/:�.�8(}�����h7Q�ئ���,>��"Y�&l��D`-af'����pG֌]r�W�f�V+��72�:Fр�N�mL+�~��nE�T(�C|�tq�?|)�Rڸ��ܲXvJ��1�=Z(,ܷ��X�`�f�����M�fz�n�KZ*�V�ֻc�T=ذSB5�����g{�8/����� ��)x&����H���s���LN�ZռO8�T�(G:��gcǝ��(�6O��֢�6������7*TW8��$K��j,
?O�R��{�0��AA���=Qo!!m�0y�g0X��IKݶ��Ėq��"��AED��F��������Hq�1{~�����$b�In�
�*�[���p��w��?����7,���'���,�n�hD��Ѿ͉	�/<-��Aw���OL���!���QP���ON�������Z-�R\���|�	 �x�x��ǖ�+Dk�]@�4!��Ze�h�E	�����T�~k�C?��V��vzd�Ό�'w��i�^�� ��M{a=*]5��p���3_K7!~��2���5���ȹ���0��U��T�b���s܆���k�<�� טq�LP0��J5{2��\������ig#-����v(����"#��|��=D�
��3Y��}���`��y��)㬃���#��:lҾs]�0j�=��TW��W�'u�RX�D%��p�ː~���B����Fk��s��7�)�2{�-��$[U����uHU?�����H�s^k�q����.�٬���~�xl[h��c�q%�{i���������Qy���&��亐���J�9	'Ei���:�Tv�"�A�`�V2.eq+�'f�U�,��gf���w+cH@�wa��7eb���h�������H��XO z�C�{��:筀��V-ނP57��>�Y�]���U�x$�������}�BA.��,��í��~���eC�����-�ӣ&�5�Q��4\^�[`+��E���xq~e�,�p�8���=/�*]aX�����6�*8���MZ���Z�=�b+���z�T禜;���.���3��$����N��[��\���z{J+#�z&�/�OE�,�fX�v ��^�h[���s��f����@#�BYW����/�õ	�F��+��!�~\Uٜ�8xm!C/�j�y����Yj	����U�GV��6�S������nL�t�qg��}��#�P�>�"�������En2W�"�?�fy=ֆ�8�陶�i�&eah(�(�OF�X�����G��i��a5-���s�@�BZlq���f��Hn�ܹ��.I�MNY�^����pc2��*��`M�- _�qy�ey���!��4�l@�\�u|p��P�ti[`o�;��]۪�¥v���^?���q�H��*�ne�5Y�%b�яꘃ� �U�&|@Α��.�V����W�&*�������`Ĝxs��E�,�x/�&���pw ��(���ϴ�_�gx\������P�R�g���x��+��B��P���D>Z��5G&Ƥ �m����lF�%�
Yq���IC�4,ꃃL�#K.g��2x�菻�pv,J���g�T�8���>&�k��;/��\�� 4�'a��2�p�(tsQ�o�_��G��p?4��g41O��`,��[۠�e��F�F�㪡�����Eǻ �}��%����ȴ�,���Ց,��5�;sil��D�P��3p��b��6���juB��E��=��'��/����� �?�7q֑7��s�� ^�nq��у������?|	�|�]UYf�0IT��|;/�Q� �~��X�|9��2���v�s�h���!�+t=*�a��N�*+����d����$�� �z�����������	��jA�ck�ɱK���#^p�sa4�k�/�_��1�~�+�
%���wM�:��ū�L�E�p�
�$��V��U57�.eT���a䖇t���~uQ�ҩ�U%�Qa`����'��(�Vx�6�(t�G�g�
����nf�fj�Wa�kA�HP�]�N���F��g��a�H@,�f(Ll'^���u{u˞=2���z�'�o6��zゔ��֔U��1G�Mj�tSx�q,�߀�c5wU|�_�\�SI� �i]LM���_-�����fv��x����4+� ���dy�����k��qy�P��@����`�,LK=$"�R�޿%S��9�I��"���B'l�1^��(�<������7K�� ۀ%�N� +��n�~w���2���P�Q�w��dU��j�D�k�r�3�&>���ht����iŲ~�y���L�o�~�En讇�P�^�W:T]�ػEaV���gz;f�b1YL�|��M�h ����x���X2�Plʦ]�J�^�2��u�1i���V�^��q
x�|�b<�ĵ,�\
�M�1(�yʨ�����z�O�G6�/Aib��1��a��Q>�,�����.Ll�J���`)P: >���F;ɀC�%��i��8UD�,��8��Гl�na���7�4N���|4��jg�?�=�2�<��s.��*�� K��}9���*�ȕĺ*#�3�R�@q�7fNǤ}�����e,<���),��/S��6�htꗷ{%y��׏���;�b���![̰��qșZ�4J���o�7�v�ߎ�m����dr���kG�GT7�(�B�h/�M-'��!(�UߢS��ڹ���0@?��U�X����C��:ʎ�߀�� b	5?Sl���ݡ2��N��M폫�p��m��M63�|e��� 0��~�뵧��V8��ҹ�B��v闲N��1��1�w�$�}ze@ã̃p6��{�"4jq�j��ŉw�[�i��7+!!���OU�Y�!x!7g��Z�r�T��rx�S^�f���_F�Dᴰ��&=�
����z)��o��"��c�S����q���\���$��_y����˿t�|ڸ÷���z�.�L�Lب�r�2G���Mõ�X�7]��s���5?�Ҽ�9�q¡6-�x�z|Z��a��[�⬺$Ը$I1MܢK�d�e�3��y�N��GC��x��U�٧k��	e�:|��=S���@QJˇ���������N�{�xs�yWb��]���ꎅ͘���
�����Uxˬ>/Y��s�^�Dp%��	�hDZh'�S�W�4|���0n2�+��ƈnb�7��r�w]jlB�r�+.�D"���i��d�>�dqn9��p �Mt:-t
�\��pD4Z�b{	y�"��$�벹�<Գ�;@��q:9�A��~F�{$s��tJx���nn��!)A�&��=Y������"�������5ۜ��X��΋r��{_�g#�d>	41I;�m���Z��֫$%��00��X2cA_� ��_�}-����=�4W�i��ȍ<�_:��K? ���.�%�5j�(YP@�Z�q���C�ÉǛ�Jm)�\N���| ���zt?�z�,\�ŕ����r��<m��\��K
*5P�M��� �"F3@܁����h����h;��.]%������
���q;��wQ��âa:x/.f�5�I�Di&U{�1c��sg<Y��Ŗ�Y�&�-XQ�K/�.�0ϗ�~j}��a���YY����H�8� h��8N�!�Y*�j�"
mPbm�G0Z��ı0%�eN)��0��t�v���)R��sO�׼K��}z��(��R��d�d��^��1 b�.2¶9Dg��X�\�t��>� ���=M�fGH����\J.j�c�B]����6�)�c��y�o�ĳ����A��n�8��<�{��=LIt��n�j�a1�5��龮�uٮ�Rad&/G��vC��gCE��L��s��,N:���c�]�[�_����M�N�����Hq�;i�2�#���ؕ�%��~��]�����uTo*����%K�/Wgp+��3v������ ��j���N^_|Ra0�6��e�����.z�m��x��r]?��o�W�)}���K�2
��
�����2P	�׆��,��dd�B�JZ��=U�i�� ����Mw�5���[�G��G�Q"Ӏ���bǴј�=Q��|G��F�.M�&�h����*ĝs% Ð�����]�G��4!�LK�A�����+/��r3fj:�%�; {Y���]�Z���k!��������g�9k�� )Esn�Uz�8��ܭf��qĥ����3O'W�΢=Y��b�e3>y=!g���y��5���kR���(�I�[�6�V3"���v
��T�4	�]a�Ly�[��͜dI©g�Ɨ��[��B�hE�ӎ �r�����9]'�����-��!W֌炕�xāЯ����"N}��7Of�+�k���e�F���<Mc�d���a Ǭ�ٜ6e@�,ς��L�p~M4U�n��c�-����y%�r�j_6_�����&~[0� �C�4�po�@�H�뜠-��7���0�<�E�����b
O�wdqBie�d�6�0wv)��P⏾tcũ�;�Z�$��<����e�k��O�"֩V��m�@X@�Q�}Х#
��<]�u�7�J%\�XH�LՄП��ݚ����4���d����pvB�,��l��{nw8�,����y�RQ��:��L����{/���{������P_�C�Bx!94�+�;�8f��B�I������ڹ�*(4�����3/���D%�5}���oþM���E;~!��K�A�֞����n�>�P#�bcz!}q���X��E����3R�H~w_��z4�0���z�\8��@��`��)�sJc_Q�F@C��pc����:sg��˴~F ��#B��G��Ff'�zO�ho���}��Cg�k{t�"��Wr����'�^o"�B����ӜXz�duZc�Ǣ�vJ��,���m\m,3{0mS6�2Y`q��3�ï�pQ3Y��4Wp �}�8���$�����cݠ�_���	�F��9���2�*o?�c'4p_Zԋ��8ߗ�P����T���Qa���?�ա�j-H�f��30U�5��L��0YN��/WG Q�Y�q�xU�l�Y�L]1֊�|���|7�����NU�b�>>�S��8;�a1%��-A6��W�`)FfOf ��X��u�\�Y�AEb�,�uy*�P� ��,tw͝�,�Ӿ��ӈn�֦��徭,U4P�j,Ef :�Ƣ�m~��e��$}�$�bq�/'�?"@+�g����`��b�P�������x;��^�'T8d=9�M�%_��ǒ*k����yC-%�0s��
�����4ڐ�+���9PQ�:7��V^:$��&豌ט�.3]i�`	Y27H�6��Fʝ؞��6��(t���hTê��^5�|��`��!1�f,���ꎶ���c��a.�L�k׺*��u Q����F�gyw\D���-p���B�X�|�- ��6�'����o<j�j
iaѝ/����Vש{31�鲌��|�^��=0%B��(Esڬ����f��k4���8k��)�#d$�`?���PأzU�u�n�� ���4�?�>K�b�߱T.W��(�Ի]�p,M��j>�[�"7T�iz���B�rz-y��_ ��Z�c��>�Q�齿�b�&[��U�%���a�����ba�+�����H09����-�Y����3�O Cw$�cY�N�of��1[�Hk"|hw�@��\3&�W
�J 5��4�N�x��2`�
����a]�/3�ES�m����b�����m1]6�y�H��M��_m񫽅?ꑥ��g��m��?�>��Wsl�;��
��'�*�@�����f�%�\UW�o�HS��'�E3���|Uk���X�\1r�L&��E��k����h+�-����fB����z��B�,�4#���P�v`�����kK2 �b����2E,*z� QO�i!�&�>�.���sX��قН�#��Y(y�Ӿ�.���.<oG�D��R5�&�}���m�
���%���w�;Y�C�[�6n�"/���+��x�-�uP��>}����	������|����w�[�d��N�Ǜb��q��QD;����p)�4������yux7az�/��$�^yQbF5Z�)��C�G0�����B@�YOM �D�GI���?�,�cտ�J�ǀ���b���E���^���t̟�0���D�h\���-���z��I����r��@�'R��6�_�5T^,�4��"{����em�������Գ>T̛���1�nL��5��HItB`�Zj͍�J��tܭ�4�eG��*LZn&�v�W���?�JS%�:�ٟ&1�6�Եj�fEB(�Ƚl���u�}oK��:�{Ci{�H��O3n��_��M��y���8IMk�eu�R4��1zI����w�����*ڀ8D��u:�����Y�I�J��SM
�P(M��MY?�
~pD�ǔw6G��J�u�5*�f�Mӳ ��W
���k
财�쮢�DY��7H}.�PQR�*�r�2gQ��Z̺�h����$[GASM()���ْ�K��ƽ�6���2H,�&��»��%y��a�������nXs�A���[�V���+�RKN����io�,�ף���݀��=K�R���N(p��%����|�߀�R�؃:)b��H��es��<����7��<��j@�!�p�H&>>$�ЌI|u���?۲AV+�sn����hh!�g�	N��;w�ׂ���Y���e3t\�Gy��}�E	� 6|
��$�4� ���)m�L�5�̴�ӖC��P�����gh��`8��%�T�����|�����y�=�"gI[�Q�Ń�gy�����@�U�h�>@�z,/YoU�{���t�j'�<m�&B{��w+[���hq*��'���H��t����S�o���}ts�*J��e�%:�(�bYO����/:XV�au��u���DQ�3>hKh�U���Y5�Y�<vr2���+m��-�n[7� n�kk�%]���� J��{�$C��~\E`B�')?�������Y+�2g��yQ�)H���G�mi��%V��:��_j@Ǜ�C��wҢ3�K�]��KY�Z���a\B83��B�F#�r�崩�IkF��Զ"	��|�d+��%ի�jc�hk�� X�{2M�6K�`�Y��$�1�~q��ߍV[T�J�#��E��Ӌˁ� !wx'��'eύ��=E�g�,�Sǧأ���%������{��	��M���3�h7&���%Kt5(�+*ת�����%�/��jO9�`�׸�����L��TM6����I
�������:�d��E�6
��	�« �跼�����@@oy��z��ibk5x��}<aO�OY0�X����\�?~)<�Dd`�e��``�V]+*i?�v6�G��7�z�9$�k���(Q�;��)�9�o���Q�QG(5�C��`H�Y��UjˮQ?4<s5�D�J:F�13^0
���hh�`i{�;���H�>.3��?�j%�c��?�����G�H
{��.�`:�/��wn�}|�0Cw�đn�E�e����|2���Em�0+�2yC�'�$g�#�ڸ$iE�VZ����W���t;�J?"Ԃ*�����UN{��.8
ʥ�Yr:O�N�uū�\�o3^.�Ћ��f�܆�N#B���h4��&�K�E����(U�Rn�p�yOZ����-���R�?0D�$.���>D}����g#���_�Z���2����X�^ J�t��4����<鈡�~��lM]+b��ʭ�-lW��mF�&�&Է� ;�?b�u�:�)�P���(g8��5Ÿ�6o�zAl /g��Z����ړr:]�g\�Й���h��t�߲%�X�˰G��҆g!`+�9 \�>r��mw">~�d I���"KT�M'm��;۠���5��A��]�H��Z8=���q�}K���� ��Di~a7A�WϦ�<��DW����5��;���d/��I4�Vz��L��aD��.��McGa1����ֱ��U>���'�r�kW�C��B�}$` i��w�-4}<*f{���C���j��)(DJ$��qә!�AR	EW�e\Tѥ�h��sp��VT�+��ׇ姦�>���J�)6Xd7d����Ya0ҵy��?e��ڼ�ҝ�l&<� ;�K��T�Q(E�_{��!�|)p���V���FZN1�v-�=]{���sXxr�����#�xx9�KZ�Apd����.� ��rA����/Θd����H(���%Q�lɞ�|/2i�msw�{>��ܸ.i����#�b�G퟉�LĒF��
����]�n{�a[�V��IA1��Z┲9J�$��Eh�x�τ�Ұ�!A��_��Q�l�NT�XG$J��9Ia�lI�⻭.�ݘJN����.�����Ի2�C��J�B#����r=��/ڹ&V�����'�K_�M�^FY�U��́	��^��qJ��		��6s�k61�P��̤�TF0.�XǦ��۩q�U������l��U�W����wrO��),8E�ܳ���H�Z�����3h�Ѻ�'ܲշ�>��69%+V��ڵ	+J�gBe:w��32�5˚��m�ktSm�*O�r[����՘��T��Ѩ
������~�<�讅�4�k�gS^�~)E����]�@;���ٽ�~��>Y�C��o^E�O�B�ߴz>�������}�iT��5�T�\a�D��k���B�5�`�U?�
���O��q��E�t���+� ?˻F��g���n��Iq;U_�'�������I~a��f���"�vWKpVD�]�eC��7��{T=a�V�z�IB������B�Ģ��9���j�	��?��j����ߛ�S���H�!��0�2w�Q�ZO�u�+�q����S��M8Hb)�|Pn3�)���'�z7��k�X���5Q	�{N�È�{y4kq�{�I��$��e&; L@�B��*6�[���p10�z���m���G�w@ɋ+�����C�V�E_�����Ȥ�W����c5�
+ćw�����d��칉��3�U�r�4�5���7�0Q�FSs0-���a��M�L�|���Յ��F `�\/q�J�L�E�Iv$B�S%�����^?��x?7�(F#���&�[�a��f��P�l�HJ��N��9�}�C�*�|��/�o.@A�̥�al�8�oX�����U�[���M�Ƭ�&Ӈ�d������-�"+(*���|.f�k������_z.�?�ͨh�|�{�~�t���H{L&��>\M��;A�Y[�ǣD������~s$v6��R��Kn��)���'�{�?-�X�2�	�>��ԃ�rv�L�&�����ڎCiZ�m��a��Ҹ73&a�+*�40�k�0�YQ̑W��<z��'�Q� X_�<����5����A_�;�HȶVW�	T����,�|�;h�:������}�w����!���_�B��(���<��f���룻pt�����ᖀ�&��9g��	�-�o9m�KiF���h.c�2����z���h(tX{�zh���+dy TB ]�LY_ݳqTG�i�P0-_�S`�$����*�#,a����p�g]S�,]W您֛�Wf����v��~5�x#�հM�eݖ����>$��И-�%��qB���;�d=X �`M�mͷ���A�a�<����Y{�v�1A�\������ڈ�CE���T��%%G�9�2�q�m�xXzJR��dO(��a$q�0��,�E0�+�3��	��s.�j3�*�M~vT�q�f!�3���{�A�@�Z~��ɑSW ��e���;_�*��NA��@i����Cy�7z��X�����Ic/��4�ΘK��z�9���~*J�W�}wF~�J^@�U��Oݫb/eN�v\]xG�qdNg��߽a���Ɔ�7[)�h�'D,�|V3�`�2-h�^Wc"�f���x[ Կ4����b�|�M�|��c3%�vM�7&���$U��*�tY'�419D1�ʋgQ�֎��1�n����i�&	=����:3�v~d�����[\�zux�zj`�urъ��=
!��o�6772c������Y�UtW*�<��ô�]2��Gm���+�gn��[�5�s�T
��oU����ct��x�4 ]�EdhlG�C���bFm�o�皤B��{�'X�FL�l�f��𘣲h���W��ؚ^�X⯏���SV�����y4��,K�
$�f�,��� leRO����ξ��ǐ�!�œ�	�n.�e����aN]Z��	�OnH9��L�j�{囍��sK��P�8O5���#�:k�
clB)���7X�$����֕C>�F� ���17�45!*����e3QO��5��j�T��&	k�59��ǧ^d1~ү�9e6!�d"{�3��V|���HbT��ٚ��<
�n$(�G�(��Et#"�S�	x��/�	���!��e����'�h��G�!���{�j�+5�r���x��*2����ǂ��M�@����!���ߚu%�A<��ǛInOY��ɣGW�L�Ǫ�I�2��kz�.pp�8ŧs��M���*?_lƒ���B�����A�E�"�,%Y���ܑ���j�`F\�`�X0�����'(%#Ε�j���`�6)BO
}�)�BEXB�*l	��a�GI�$h%�����o�)#��	\G��c���=��e�8�	8���A�z��e!��]�23���~un�� NJG���e����@4?��gTW@��zt�ϧ�#f�MK�AD?��p�Ƴ-+�#�����_�4ӓ2g����;�W˛>�H�(��2 gR��⼑����hx�|LPy�k}�Sΐ�a�8: q���F/������/�����pSw���	�(&jj������T��oD���� ?�Ճ�J�<X�D��ó�P�a��A��ʵ���{w�_a���)p�C��]�͒{�;���(��
꨻Z�LԀ��BBG��˯����*���l�2MK�R�٢��_�M�V�)���v���*�7�q��6�0E(D�`H$F1Ap�����Ħ�̡�y��g�
<\�y`}p&�{����
�U�"��k�5�&�N�xl��B��6r�l+`9� �)����Yo����Jwj����G#j�9O�l545A�>{�t1y�9r�x����S#��#�H�E]Qw���˜-k"!ФC�S�\�����;eIbؽeb�R��9~}���WT��"�@S�01I�@ɵ�~,�A���[ OZAl��}�8O p���	�ԜlP4h>�%��L���i�--�e[f��«(}�^]��_u�3���� mg����*��5C+�����Ǝƿ�U/i�M� 1������XhQ�T4�\>��/>U.��W���Il�
�#U:g�l#F61���ϸ(l�[��b��g,?gT@���,KQ2�V��8�=j��6a�?�p����t��<���R���ꦡ��&V��"�"��f����B�B���p�C�f��L��<���\��,��$�W�J%r�� �S�%Y[�V'la�媳�@ߑ��"kW���h��[GXf>DT!x��WQ痄��8LM�(����S��]m�R}���-"B��Z+�8�N�Or^�TupJʀ�׿��T��p�k�eas�3y�t�L�r%�5󅎸�h��ΉIV���<q�yǟl����h��gh�\��	��5�K�.ɂ+ NEG!�K������ϺQ!<~i6�n�9�:=��ib�O��gԤ)b=S���]10�JJ��C�0xu�n4p���M3r���~%��KBJ�g3�9�m�ȁŜ�d�f9K��΢��w���A��'��Y��մY:�B�Ŗ{1X�]$i2�M�q���l��K9E#�`�O�bEXj��d ���I7#�J���ID^<�heH�2����-y�����ԫ�#��P�^�%l�s� 
���m����K]c�W�m P��ZC�sK�����H�y��[��I�$��C�xe�^�2�s�c���d�i��)2񥀬vb��`J��Пm�����#���/��XG۷袹�쳃�`s*����;zS���X5%��g9$�B�s�;9��_C+E��<Rj�QgR�'��叛@�/����Ć}Cm4F;4og�P}T.��k(:�#���9sw߈�D7�[��n��3:�GC��llK��h4����2�ʹ���j�w�9���f���*��d�ף:�}Mè�ء�mD��šuK3x���a�ۻ2Sp��]�-��=��&��2��x ���R�!"��P�ha��I.�j�����4��ހ	UT�a:K�'�-�G$I����Z���� �K��F�:Y���6���
�c�G��Y*��腑���MΌi�Z�AuN��.%]2���Jt�X�
C_���щ�&*���
~γ0���ד�Z;���s��<�Fr9���l:,�YMc뺕FP�&�V��i��)��X��GU�)ݭ�?
j��ΰ(h��%(G/��ک>�Y豠�Ǖ9-�@�~�B�3�!c ~G�(�����ҏ|�c�8���A�d�G��-+�sG�j��D��n����+��;6�ょk�$��C���1���<c�j�ኤ�����Ġ�f��9:R"�� �g�4�f��e�n�Bu�L6U�y_'��������E�a�3�A��H�2vd����`�AQ����&�EW��!�_��ґeM.ƣDĬ�̓O�rM*Mh����G�l/m�+4��63�H��L�$s�s���f�!��U;u�EK��x�������7�i՘[�1�P�"5Ϛu�����|t;^��F��|��osJJ Y�h"�~}�-�&Gdy|���2�S�=�����YMM9��I�}���2��xK��0�d秓Bx�����i�:�K-��]q�����hͬ��*����Uk�X�%2��Ա�0�Kc�q+X��X�r�H�L��5�*w���nUD��拴�,Ms/�8�|��A���E��p8RKa��	��������s- +x�Jk�j�zJH��ꐗ��}�'؈�:ꑁ6�E��@b���iny�Qf@�[\������%1s+Te�
��.�s�}�),�H-�����	�!xd�t���'�$[��K����P`��C2�=/�u��҆4O�Ɏ:�
�/�T1e������an¯%�xJZ��c�M�a+���o��L������3-Gr2Qʣ�`���5@�G��*9�\m��]q��B�mN����
[��g#c����(}������^��R� ���dj���K��*���;�����	����1pKd.U.3Pevo��u{S���=�׵y�e%�25��uϥMG��,����.x?��%�YIά �'�V>�r4�xh��O�q��Q*��|u� �Sr2( �ba\�_ns# ~%?f.I ���7��u�;��p1�fQ� �Lt�z��ʙc㽜K��%-�[U��R�`�N�e�g�������U����4���1p���Lw+OR�G�q�\��/=�a�?7[:T�v_}��s���F�T��e���Gz��v�}����#r(���)?�ĪjTڢd�IC�����'�b,D�,<�\tW��\������B�V��I/� ��%pY�jU&ѫ٤��8W���cyy.V���{��=%8�u��h���Pfuy�)�>7Ŕ2�%O�ߙ5��s����.�@�J��٣�OX�+���:���@Z�b�U��ɯ�V�(�98���6d�y�|�#8[g�CR�p���:�k�J`խ'�՛���{@�f�'��h��#~ۇP�v�*4��#��j��}�|��%���#�?���? uM��ь�_���d��b.�I���F�~;D$�E���r�/c�	hb��b�%8���7CG���������l(��gj�W~�r��Ă)I���"������	��e[�>�L�w��g!o����g��<	��^L�T���.\�Yk��{���!\�0���Q�t��<)$34@����p�=����&�O����y�"ˆ	�:����pO��!bN_p������4� �hAD�s9KX��Y*���ز����v�I@�B;�Q���|�m��yo�����62�x���x�u]�u"�,�7I�7e<��V�;��Ć׭F�%3�����QhҊ�����NCi֧h3u�ބ�Ajy/����y��a�m���>�����
�@�?�� 84�����ҳ)J�
s�W��	ab��v/�\n�DЏ����Q�ʸkJ`z������J��R�v&4R4�n������z�c��6!��!j>���]�{KeE�aP[��c���K{p����n��{�+>��ԓ~��/��!�d�Z1�?�Jm��Bn�$�)������h!1�xNsg�E�O�	��>d���SZ�U�v�)(t�n�F����˸��v�|��#�3�����r����8Q�\w�z��[���M:)N��DD����M��?�Y����<�҈���L�KDU!x"_�5�s��s���z�	�|�9{�~�k!�8C�o�&�X@M�'�Չ�C���S�F�� 2^���G��p%���Z�Hr-�����C��"VIlۢ���Vx��Oy�
M|���N�#�ğ�����hv���u��m�oQvQ1'�1�ǉ��H�Pc�����s�rs�L��tBıT���[i5 �݅c��k�H��Ǐ׀��2j�B�m+��ɚ��_�25I����;�w�I�Վ��,��:�S���Y��Wǆ�2�%u���8w{�~p����:�����'\��n��mC�쿬��
��P�+�]��D`�O
��Db�P\�HPT����h*��L���\�F�݅�:�m]knSX��Qo�i-��hHMD}b�c`�Bt��_���*)ͿX˘��ї��v��i�1��� j	����:�y%)�F�V��n�ry�˫��§��H6�R}冷/�d�da?3z���cn����J���3�'�����u���R�g�3
��C�#�C\��
La�ފSGe3�T��J0����W�9��ub�bFE�hJ{"��P����S��=Ꝿ��kX��o%�-Ї���翄۽�W&�`7V/O�a����<)�w1G�ᆎ��;�܄��;Ƞ���bFa�b�U"j�`R���NX�nR�v�F�A������fa�c.ʨ"<�/�-�F*�^u�Ď-_=�62��~\׍���Qk=��3~�ii��>�^��E#���
�i��3���O�W+�c�0�g]S�-.�օ�;@�O���X�a>�z
1OIf:�6�G�u:�WM1m�+����!Y�5D��'j���Ƣ������������;�������<�����OA��+0��$��!yԮ�g�Ev��e�w��t��N;e��v��������)�o������H�2
"��,j�i�	����'Y��6@C��I�d
����Mq��/t�	U�ڔ*�B3��ښ���2�dIK~�( ���z`�e�B�(
^������a�i�_�=�?J:ˁ5LH��8>����m�&�$�,�1��tA�����F�I����0�J����t�&����K�E���eku�ج>�!��gOV[��zD��ޓ�(]��ׯ�f���'R�Sl�3F�Lv_J"�T�wT�'�CnOE���P��(�`�u�R����u_ĺ/��Q$��A�L'�� Wk�aVc�5W��Z�7L�/N��]희8s[*����-U���Ӛ���h����e�U�N���T^9x��m�PC��݉P�P������G8��M��+��k��:j�̬�;[�e��E��	nQ?����S�;kI��WV�LQ��l>)s5�8&_�n锅#H�!sg���gy[ڵ�k������ ����'8e'֒���?���}��qГ04( "�7�edV�+�7����� �]!d� �Gu��Ϩ��O��GR�����p��6
���lkB3�2�1)z�(yNJ������ G C�*�F�Z�@^�3J[~���[�������Y,q P���j���f���TA����,�X�\i��]*���i�u�"�g������>f��-������,5ⰾ��D�<�Ɯc��"i�W�}I�>�-�F9�%^����0����ҹ D(:�A�M�/����a��PJ,��B{��4N����1�Hb��
7P��͞I�|���a3�y1�K���/)>;mӹ����5�@��m�H}�{�&�Ci��"���Bq�D�,�#�;���xa��ӴQ��o�"�M��-`Gw��8׾Kft�����҂*�l����*�����Fr�Y�e����OIj�B��)dHs�U��n*���S/1��/ju����
w�^r⧑
���NYc�#+���E�,�6�+Ghf��3��:3�2�2尔 8�PQx�Y_!~��G^B�}V�G�����t<G�1����� �@���k0r������U�#��E�$s��"���$v���rY[E���!����8�Q���; @��WS��}�?'��ڒǦ�\��LH$��
X��D9���4 {^L���{�1�.�S����N�:�@b$�,1�v.������r�E� F���D���j��x.I���On���*�G�N�W��r���t���@�Z��xqB���3�,��<�!�r.��~���jf�nK�֡�5��Qm����<h��� y���/ �?2+��DW�g��UDՅ�r���g��8�_ c��Z��|��){����"�$-W@��A�q�u%��,b��%>�5r�M�:��������g��N��~i��X�{�����B���Ŏ�<س>��Y��Ć�pip�<�p���*-���{��ڨ�v��]����D�1k�P	dB�����$U�= ��'�j�S�#�5r��J<e�	q���JS��9�G���:z;9���_4d�R��}x�bu����Lp6��Q�$�dv�v��c	�i���]��Y�-0n�Jc�$���q$Oc���>����Ȼ���{��Sk���`�aƬ����%T|]�=�`��>��c*}y	��f"�A��.G�eh�N�7z���)������ ����o����U�m�CC��M�*ޅ_Ȭ�Z_2��s8��&�1�grv�	We�J�(޹�\4�9��%�`�틥4�$SU��+�e�\�iP��.���B������Ϭ �ʾ�x��
�KΡ�DF��~�8���v��Re_;�(�.�>�A�R���)���C	Y�Y���*��Y��� A��H�;?L6�4e����gFi�*��!R\˴�aH�HcoR�@1���÷��a!R-%�3������J]�����G����׉m�7���Ɵ�2-�mFkT"�Z�J�Q�
*S����j V�]��-�h������}XM���V~�r5�]�;����3�;�E�"�'���1;/n�HҀ�E����t6���s����2�7�'Po�dAb���&���{A�amS�����/�a;
h�qa�"N�aW7ੑ�l�w��y���b�NU�C{٣Ar��ʷ���0���l/��MF�ޚ�����1�P��k�r�Ѧ�m�0�aX;ɇ��`��y�2�T�����ؐ��Z�x��B����{AB���y��99(B��ȯ�Ţ���w��`��u�Ev2�l��kY���K���g��������L�?�p�*�i.д��i
5�����B�-���^ڢ�	�ǜx�B�*)s�>�l#v?G�mk���t�LgWRc*:��r� 9�c:VJ�*[ηa}6R�Ώ��ߛ��Ό���8�v�K���;���U�
��^�RT���1S�Ot8GU=s������|i1�5"9����2*�v��ۅM5ہ��!S���4�	�ݶ)�Nz��#�B�5��~Y�#G��.OG5w��H���I�����9x��4M3o�=|�U[�b|lX$ükL}k0W��]A�� ��s�C���VuT��~d���w1��{��DT�2�͗�_��و�~׳�ЛK�H�s��P���c�%��{9�ѝ���zT�1Ґ��d�S�ٵ�b��Z<�9�&h����)39^8���C������P=��8�E�z�����ܮtՅX�)qO��
�)��u1�+5��%<���{����ue �(;:�˛�cd7q� ��J,�!���w>�!ն#���=��/ߎð�و"�ɽ���3C>�� �TM�����L�f��X+���x�w3Q(���+ó-x����ߒ"�엧v�La*��>?32����R������$�T�~?#�Y���R����1ۅ����2NCm}�ro�\�9rҏ�e>h��/�J��y�j�k{���B�����+_��8=!.Ek�p�s���ɖKR��.4u�W��9@��ܴ[�֋�����Z0���^�*�C^��ZW�����r�j�B!�O��:��d�29@\��!�J�7`��P��
6��2��)g(�o$���������X���[���(����ܵL�B���O|}WM���;HQ�f�S����B#�F�g_������G�d�������ܞ�2IU��Fu�1@��C�h(��w�p���6o�'̷�mb��b�R�.��wrs�-��#i��eET�,��H&��Q�\�T�$�䬳��h�9~��a�IO�[�88�ι�L���I�M��hAg#��}�ͦZ뀩��o`�92";�r�	2�z�౽�7��=(�"��,�:��r`�8���jw��b�	}i)t���9�2R����,�Z�ފ���.�lU�w��do�y�."20�邿*������R�Gxd&��h{���^�Դ[n�l��>��q��HA��@�� .�e:�s�~����mY�}0��+s�R5�n/V]�.���h�akڀ(f;�|���{�
����[,b蝉ݬ���'2=�t�VxP=͹ˡ�ю�jI����G&!���1�&�HŅ\1m��:��5Z�)��5^�n�4d�`��
M�ǭd���K��f'��)��ֺ��Rs� Ϙ�1�X`[vJJp*zW�NSY�fn=��~��d����ES�$[����+o�����B����2�Aß�<Y��Ӝ��K�k�_���h PmO59\�kyv8�yQ�j�g��A��c�s��-�v@��Ec�C��4�Q����]��*Բ����7֥M�\�!��+�F��9��TWd�����SG2���aǼlv|�U���E�~���M���0�K���K��Eb7*$��)}܇��d�
3�҉�m��n>q�}�f	^����2W�*M�<+ ���@Y���+x��^u����xˌ���'��#�������Y?�l�TU�3ٓ��?�B�63`����ȒƦ�@�2����X��.���K���������R:è���R@��gc��6��Q����\��lߜ�T~-딝�s�Y�)�bW���d�[7��������4�}�r��q�k}�sC�}��<�ѺH����z 7籩�2��O�Ji�[���(�6����������)O��N,ڧ���3f����D�#Ʈ��cDn������t�uHӜ27���������r�|�I��X���	al�q������ Ą�0����""���񨤌�"�Tx��� ��yy��%�B��@�Z|�����y���@ϊ�ޥ^G��r�v��D��}9�cE#	[���hw��w8}8��<2�޺w�J�M�}1�Hӎ�n+�{� �O��x������ǯbJ�3��E&�����
T鉾�v�?_{��k�1l=+�j{�F�cס�T����=0=��`-*}gU��oFOw՚x�;���zmCA�5r ���	6=fT(���A�[�SX����շ�^VS�kSl�XrkfZh� 
��UQ_zo�c�?W�d�����VI��\�;#���Ӝ5^1X��Z�'&��>�{+*�p���	����uĄ����ኬ����2(�5�����f \F�%|���d��Ԩ�$��O^,�Y	�y�hп�HQ�]tr���H�C,*CFX��[p*��!P&V3zI,����u�k��'����=MrZ��A��w�+>�/�R�n������y�?�Y� 	;��RS���ݓ��)�5���D�a�H����D�?�UXNׂP_��GHN�L��� Q-��e��D��0S ���I�]��Ɯ�1��ůJO�#㈣q��
�x�����l�2�F��CAT ��J�"��q�32�k}�8q����SPvX�m#�9;F��z�N9��*�Z��4C�ê'��=����ca�<���/���������X�>�Tt7uhy�C򬳔9�K���F��"!��۷	�'`_�4dy���|�2i��Ek_�Î��z��ؿ���{;EV$�o,��YS�Lu�e����ϯ��[��>�Z����8��c��GC�G#��ړ�PN���#h9V���|7�ު�f�3_���Х��t�"�W �3���hŀJ�%@�l;�=�P����%D<��!uY�pU�Q40��tj���f�T.0��јx\�Ɏg|�TL7�AAz?��h(�Le��
?��"�� �A9�8��?x/��?���strI�9M���,����/*����Q�y�Ԏ�1��0��t�I�z�ɍ.61����ttx7��̉%j��MMAh��S.����e�d��!N�����$��l7��5� ʱ������`o�O�K@Bhew�����^�M��fOQ�N������J#M���𕃌�*�ݒ�:*X�{�[Ա�^�/X��]a�Ci!����q6����N�R\�&6Su%B��!�<w��ħE�Y��Z�nՋ�k��m�^k�C����m:����r��?p2���Iн��@+EI1��V���	����`����*x��m��̻J��D%y����qb�حmG����5�u}�*5�yjɝ��%�摱���E뿰��o�u5��u��rfɄ��������!� Y�W�����K�|��cj�OzU��f��֐G=I5���ZG�6e�n�vK�,�l56�u"5���E�}a��PI;��Z�띯��k)!K�3�<��^H�wɯ4�?�z� B˩�|���FeJ�djm1q4 �1�G'�,�"3����*�n�� ���!�����b8���bӇ������K���p����H$��b�)T2��cz/7[Վ��?�`�|lp�6tߣ�����Ԍ�'�E��J��n�Eƺry@�	��
�N~>�$H'�W������`AQ��M)�&=�D	�44����ך��eĲu}��B(Z#�{�GU�a�}��=�bqA��1�Df��"Kư���cW�S,c��hN�I��r�H��U��V�88���r0�z+�o�@���	���ɖ>�s�H��, ��Na�0�|F�.0(�~!>��T%��Y�Ν��^���
�FI��䆶�d@|�%���V�-Sl�|�S�8%�&�U��j8���H��S'��)�>���3X��h���oFrx.�Ө�&;�1�>�f���ځҙqK�O�$=K�L��:��c1�C���i$�\��OZ۞]	�y�^�(0�Q
UPμ��&:���G�e̝���H.­���H+�MR+AH�}�l�30CA4���
�1��.�R1*��,�@���^P�ME!��
�Y�j������/��]����+�xP��������'�����<�$���q}�.�Ȇ?)������4�֤Q���z��xV��.�]6L�2�"�+�}lk�4�%P�=�k�f�qǑb�v�}�P�K�K\�h���-4\��c>��FE[�е��3�*��pn��0\_�гߒk�j-}]hsW��������U,��v&�V�W�o�{r��F��-.<��^P8I���J@^sf��2��I���H9<��ml<1��t���a�WIK	[��?�oNV$���zi^w�<�ͼ�3��Vs����h��ڄ2����\k��=���Q�|(��P�3��)/����+g��@��>�\#EdK�7�
�=* �iX�ms����VN�����Φ:��w��+`E1w��f�YR�>*��?^h����"���r) ����t @D��z�57��]�����@7�:���	�3��\'�(:VQEڭ��[�<n�3헲K$r�W$x:�?�]����\m�.�ą��ff�{�.���hp|��D���X/�@�=OIH����W�%֟��*�a����h��U�~�-��ቤ���f���zY��/]�/��d�[�,�	0��׷�������p2����)�zp�[��rwm��˔����`m k �c|�i�`5��c_DǨ�
�F�����p���6�
��y���0$x�}L5L�>x5"{&&��>U��T���S1ƫ��~S�ܺHw����>	Z\�q�R>�+��(B�V�ubGg�ܺA�,��w�!3 �m��qY�C	7���L�p݇�ɉ��,#f�|~>�YDiJ_�Q�/V,����,I�V譨����k5�t����q>W��g��ݑ��M�|��	f�[rA���|��S+�t����Lj��)�W̷��|������Tb��Þ��ڟ��*-jͮ�
���=�������K�1�>k�!ZU���z<����q�1���?��iD{{6j�=t)�_��y<a�	� E?���a�F+u�ň��A�_���d>����ϱ��H�d;�-�ZX
D�r���Y�zRE	� F$[�5�W��ݏ˺���*�<u�6�Ԑ-n�Z�\�%p���<��=���qU�?;)��f�\�S7f"��:����tM|��I7a�A΂!&2ɒ�)M5�d}�%S7��6����t�%�� 4*��>que�_�6Q0c?ɚ4���d�B��KY۶�xx*`%� Z�コǺG
�:��>+k�^i��#�p����@��̜�m���Q��IY$�;�r���c�C^�¦�Z���uS�& ��6�6̕����Y�bT��,�^��v�1�Q^���B" @T}qT�Z[�M�P���j!��4���s�hT�Ҡ�/�*f6�6&SnW4`�����Z��ڡᡁ��ٲQY�Ź�E���W��>p�W,'+���]��ׅG��4���|�*�pc�.�5>��VKV�4?o0a�"p��=�G�O�ڠ)٢�:�?���k�e��(ou�ǖ4P^�R���X�ݕ�?�i�,�u�v+��C��]/ϰ���u�����j����k5�T��6_��k*�%ډ���|������ӣ�`��&�~�~t��Lg��x�E6ʜ��9�� ��V��@��� ����x	�?���^v��ϐ#�i�Q^~0���g)î��p"�zoH�HFH�`o 4�Y%W#4F��D�ώ3�y=�՞gEr��±��h��`��p4���/yR�#�R�����ʊs-a!��Ve��?�<��t.��	l�>����R���?L�OΑ�i��ǚ8�e�!����*ɻ@�.�{S��Ô�ֻ�� WK7āo�A�v��72��� \Ϥ=T�]>\�!�]�k���D�^f.\�V��=��1�A6XR(�ŖW�}Eu�����^���AW�	��/< g/O�V��M.ܲ��2\��PVp����9Q6��f����O<�c#x�{�k���� ����e��7�\�=���1�L[!��KQ��{'��w�\��N?,���^#�Ԯt��})��vWx}�۶�s����~De�Mh_r�7y$�|�j	�{� �}�`�g"m�I��"�@�Ǩ�x"
��]v(��k�Z�٠M�y-F��R�!�]�ޅ���z�@W������J�C��Z��"8��P��d��c�6��e��kEo���yJJ�<ȇM���o Ǜý�g��y���/(���C/}j(6�v��D�򱆄ߣ'~S�ta1_N+W�3$[��Ҟ^Fq�x������S:�8Ϣ���Χ� e"�C��ϵ��}��CSl�U�Z����&����3�3t���72�ˬ��x;�����ġ�p藆�ʫ��o1���l£!��G���f �=v<�^mt�7?b^Z�V��SD/��`[N�}\o��������d4���	�p��� ����G{t�$ђ
�68Tʅ��4�p�@N\�0Y#��Y�9ٿqz��?�ǒ�k��$���^�&[��=�=΋�]�@k�s��a ��B�*���ԅ�,+��:XF6��~��n����!m$=HA��;����E�`g~4Ċ���*�F��w�1>���P@	���:���ߨ��3���Ͳs1��2��p�[S��i��el_I�=�%�4D�c�Y��\ �%�9!��@|1�|��_0J�JH�g���^2�啍#����(��� ���w�'�g�J.o��&d+��閞E#坲�Ƚ�{����D���7Β�����=K�=��/�XyV)����O���]�1���������
�ൺv�?��߈��1x�[��aNK��`8KՌ_{�6(�@ܚ�T���N_N(��٦�;Q>#�׮1�G��ۢX���T_t���w�`V��d�TKJp�Ri�_T
��x�α���73���zLPq�7�e���	�v��� �	�
��}���9}U�M��$����?!L���%��P�7���r����1��������fכ���Y�!I��#���?`+c$�����2�`&�Twn=�ܗ���	aNeQF��%(��$�\W�T�e�a�V�4%kI&0��{v� ���`��!M'u��ݥala��ZM/>9B�x4��gn�J��K�8���sѻ$�)�T������X�;&��������X�aߊ��'�Ħ�h��1[Mw�;�A�-�^���?����h����v�歯��ͷ��1������|��W�9,�VT*���)}y8k�H0q2��m_��󘠲�����	�))�*� y3��r�:� �W�dĘw���,&��H�<���s\jWqS�BG9��tN��5��X��6	$�`��*m&��l_��/�.ڠ'�9�Q1�d��ԁ��pG��ca����،�����j(�D���=���/��8����S�}���������	��u���)`G�LW,Q��m7�ˋ���:����A����
q��G�ૅzA��h^9H�*3%$%0V�S��q�S`�V��öb�s��jcH�����~�5��(fI�$�:FOKA��zv����aN6-<���[u��P�aQ�Ntٛ��H��F��i�Rc�(K�OC�S�"�(B�Fe����d�_?���I2�^!ƋY�ajΏI���љę¸�8m�~�6c�E]�V4���0O��_�+��y�Flȯ)�4���"�"B9qO��ڋ;��t�㖚r���DEp�W��ã�h�\�X��EN��jo�~�c�&6�������H�ʬ�TM_/7{�5��߼��#�X��V7_J�m�t��֞��~M+Î�=�}��=��ּ��U�6�o�w0�J������r��p�a�)�81 ,�Ţ���M,1Gzt1�AF�^���s��P��ME t٣9ZV
ld���c�MJ�04�q����b���(���GsTX ���F�zb�	Y���%�j�E)f>]�;�h�jԉ���5����\cᓭ�k8&o�J���y����:9'�Z�y.�3��!��؍_�c_�ći	 l��9W��2v�
�q9�����h�A���"Pb���X�lAClu������§�j����xN��!�)@�#�(j��vx�O�H���ZeC�M��1��U�i�rJ�h��N��1a�1Uö	'lL,/7z0ni���=����}G�<8V��'I9r]���oT��&�J�:nS��T�`��s�{"[�?��q)��*�ۊq�J��e챓;�j��^&3,��>��ڻ�\��)�K��kԞ�G�)E��+�sGM�@�tFL����u�A�,,��4HmH�6�՗��H����ǵ���G�W`��F	�][cmԢ!OT��R>�Л��VU�x�: 8�3Д����� �&�La��/5��$�yfUF�:7-\��fuh�e�J�r�Y]QmWih�]�]�#�+��r��GbrE�u�{ʱ�}�%5��me�ưҦ���T�M���0�j�U���ղ�`,��Nb�3�M,�
e��*��� *�I�v�T�ة�!�zb˹�v����o�����\��׽qa�Y%���
Ho��	�Em�.~V?�����B�8с��r���o���:�'�Ȉ�6)DS��{NRx�D^�`]D��J�1�$�?�Y͸Ѿ ����R@}�d�Q���]O}?��O�Қ�.n����l�n�`p���D��f����Є&�����9�p>���;����wQ����ӽ��OO�B�S�\���BW��Z,K��nf��/i�F�Vv��t)�n�fM!���GPz�0c�d��)���bMx��)�p
��[���a���[����
���XsS�'�Pչae�]+q��'Lt�H��Y|G��5��U���z���v^2���Im�֬�|���>z G�v�Jd���w��ra�$l¿X��§{���^�,�pF�
����2M�` R����ɳ�1_x�h���S(����ϊ\{!�mU��5�Cj��{�����!`�;-��B8���Wj��I�}D��HG�ݢ{���>A��0�u�@P6�Rj*�{���n�%��S�*O���n�wI
�V��(�s&�v=�-�q#t״f
?�*�RD�tc/��o��#1�x�����B�h��$=Ϝ��X�,���?����F�-T��E�ܼ��+��L����w���}S1|��E���TxZ�衻�u=$9ع�*i4�eD<�D=T���	{6��!�@EN�����:.��\�]�ֳ��(��{�Q�%Lz����rF؊g�B�-�/���l��e�.��
d=3-�~l�ΰv���u�Yu���+���ԩ���|۝�'�֐��~B��|Ur�-�a�)i cE�3ֲ���m:�n�Nw#>3mܹ�gC�އ+)�yPSF\�;F	���gb<M�|��T�^G����ЃT��No+y���pC_;���W~IN
���\ᐮ-�ad��^໭ ��_Ev��C��L�r�Ǧ̆:{l��VUh�$���v~z�o
*U�@������䋡�o�#AOnY�-k2��T^����9����^�h�R
Y��to��c����>C��3�;����}<ab��am.�(�Yb�|�	��	B��Ĵ�T�7������/a �:�9M�W2������DUk��W �B�� =�׼n�\"���,u.�ԃ]�.�����(���_с�p��h�&6)G&($��ƄDRܐG�C��{���檤OD��Yn�|��x�������-�C\B��Pq�٥��in*<�^� ���H<�XX�|Z��G����t�� ��O���x��䥋�鈜�����%����$�r��\�!N�ҭ�)��:2�(�UD�wə-E��S�,a9��EX/l_�?�ٓ�z�v[ �,L�Z��D�A_���	e$i��r9��5�n�KSP����	�.'����Vu2L۞1��0�:�]Rđ�t<��%? Z�g�m�����?Ǻ.D�$�]�G)5F���&�/��i,��J�1������v5��F��`��'!���p�@v@����+�/�«h^.�᰸< Vb8�U�v0Ñ�_0�?��`HZ鐊�5��倏���RE�5�=&T�`���-Ҍ��WqN���O���Q��=�u�U�!�^-�ѻ4;�S�ٱ��(��Mo���R�ٲ��W%�wޞ1o]kŏ9����뛭)S�
y����	
DoI�b1�@�y��,H��}�)dQ$�a�Z�+�~Wְ}�9%���}���S'��;3LPp�.�$#A�_�}
V!��i�v�2�*],�XK?r���TE�.#��M�6ȕ\�y��~H�	zG�XRΆ�۩�oT`̑R��R#M|��U��`����*���z/�J�_��@�~Q�q�	+���W��,�c)�R���6mw��|p5�1�n��(6�$.r����Y���K��
�j��⏦P�x��QaE���B����5���
�[��������CWjWEdv��r��k�]��<��]�9�r��Z�AR^/�B�C�B,��
e`�B��p|��Y�� �*U�X%�F�ǿE=8���кȯ�*�����d��a�GKo?v�=KB&7o�hm2�����=yB�%[B��Єخ�k:��/��zJ���A$@;��u�X�	��G��-@���}�=�l�>	H��w���̳��ĝѺ�,�>��zy��c$i�<���_d)�������"q� A��&��� ?>[
d>�C�2b{a�P����I��U�r��h�u����B�=�I?�Ymx2T�vyZ���e�2��^�!�����)wr�+�v�v��!SG���L:M�B��6���Q���=/�q٬*�r^<|I��|-���Uم¤T��K+��mL��|
�W>�'��c�ny���u�a���2��1r �M)�G��S�M1��Vbk���@��fK��-��W�Y;I��έĳ��gШI?�9!�*®����^J��Pu	�08hVn�G��*�K� n'�h.���ę;	z�A �՝$�����Mt�vzu0wt�M��*)�,e\��EE��	9����NGgS���i&�
��y�{ЍW��d}	���:4�����[�*�@�e�z�EԶ�^�3yp"Dp �ŝ�r�eL�ܧ;�� z:'��̨�?��6CJ_TBҸ�;�g���/��:xBPF����C�Oޖ'�8�N�}�7������I�U8,�WZ��{��p¥�2�M��O���on�̃c��M��gw6,c�j�Zóz�<���K�Q�-&yrJ�	O�3���vKT~�L����zZT=W�x�vB�~��'�D�n��p���&� �����J8�ژ�bJ�_�β���,�izq5����1���k�f6���E����L�8	�D���Ka4�M��2�!l��`��s8S�ɤbƂ��Bbr��,(�v���א#��S�?�,S!��q�0 �m���v���"�=ܧ���aa<��b��a��?L��5S5:A���p���"��)�M�9�vQ��b:�n��J�5E+��>�><���^�$��X��Pe"_
C?7�i�o�p1c�9i0�7�#� ���l��30WM}PG����D"A6�ݫD/���4�J�$؞E	���O�I��HC�p1�l92�N�E>K#�o�qX@�-��/�^v�<��_b%�p~���ࢀ�.!�#p^N�**�\d�����K�B������s���!@'E�a�it���9`n�Y.X2�s\����|FDpHi�z�c�V��A�C�JNC�R�aR�EJG�3�*K���^dЮ��4Su�1�`��3�Ka���s����G)�IIA���I&��}��^c�w�?*9ؒU-�n�0[8ǥ>��#�������@<GE�x���F߁n�3{m{Sc����Yn�℡_;E�Z���R��Od_v��Lz���J{����ܪ}�6{a��A��a�%�v��v.2��1�\���»�
Qd���{/P�uk���PX���z��o��[�[�b��,ҳ�����5-@\��0ho��Lk]��S�ٵ���"�~]Hi������z���i	O/�:(7�nd�F��&+3PJ�,��C�y��ۚ�`�S���;qB�UY|-�3��&�����p��Rf��r�w��֋D����9#�i�M�A�#�!ǘB��ۨ��}B'�H��T�\��������**��(�F�sv
�n!�<<wz��@��!�@�*k�"��Ǐ`���\u'~BO��mu#��.���;�O��2�7�"�aߵ(�I$��tp���gŔ�S茲�k�ڶvǽ��j�����)��5_�x���K�7R�7��^#����M�RA��j-VN^P���S�L�4�Ȝ�8��ʔ�
������G�P������A����Z��;���[i��`���O��馞�$2N >�mn먊��B��/姜��&�X�hR̴������/ML��ʷjDR���D�e�iK�9�n����G�r�h�dB���j�i�[#BM�5Zc+��v]�ı��H�˨�'i�e���V�u�{��F�
��n���Ah��
ے�������<shg(Q��dˉ@В�/݇�p��(�q���O����>Ii_	gW���6����Q׼k���޺+���'/m�G���?S��t����b�"�:��6_�.<���_��C���\�ӧ�ِ���%z+%^^׭�+�Ala��~ޯ�7ˀ-�
8L��>�"�|*�3|�x�r�#����e���lG\��:Wp s�)��DCZ)�K1��dǣ\6kd 3�l�������k�ž����%��D�E��w�~b�9ڠ¤�Pѯ�A�c�_To��^N�b��+NU&�R��rO͇͌�DQ�2L������V8:-`�� ����`3S�E����E5��5�������[AFuj��P-�ؼ���ْ�q��T|^�'�y_	@0z7��-��2�߫�_�s)������ʆq����rᎨ:Mk 7c�sW� n%���d8,{�"r�v����w���?Qq3K.�J���?�Ι�	~�I�Q]�_uE(��� <���Q.��;���T�_�;؅jm�"0��j�C@�"��[ $�~�4x��=⑌rʧ�R9��$ ��á�j�o�b�Ì�Q<1܎}���èR^�Kw*��Mְ̼�8��!faC�F���<�q|��ZN{fk����3TQ K���� �&@��U��++M�(o��^w�� dn��~c�*) ��O�Mf�컇S!
=
rl�2�*��L���'Q�M+�[�. \k��au030(;��f%x����|X�c�qfa����=�P��e���5_���yBK�27x��eb H*���a�Z0�e��V��J�D�pN�������6]�_e�k��t̯�6�w��ě#AZ���	:tF 
��T�����T���zE]��*˗�'��[ur��v�n�(?����p���h�8@�˛Zއl�� ���?7/�d}'m$���8W���b)Y�'�KOdnm�Ն����#�fL�Iִ�� Z�J�Ί7Okw]��*2c�4���D���&�6Jk��?R�ʥ�������Tx��I��H9Y����W0�r�	�mm�J�w+8�oḥ��P~��g"`����H�0S�5����0K�+��N�g�\Y�<�ח�1��Eɮ3�./��Ba����n
p�m�F�ч�GA�LZ.E���Wa�}?��C���L�83�n��Ӈ/ԅ�m��Etu�n�:��,���i��J��1vַ��Y�y�+x +j兴�&�[)���<��zy��2�?z�'n\_t8���;c��K��k{ť��E.�����M��m8�^��>�R|��5%w?���i�m�P��S;��&Lf)��٪r���@�V��+`���K8�P�%�C�E���.�P�!��:�]���^�w5�R)��c5�g���Go�ٖ���[�@Y�䷉��1?����N?��Q_�dg�6��ȃh`Y��<C�ћx����6)5@�M+�j�#tb�N�7�֐j����ln��f}��6hM���� #�&�0�I�u�HW,5
Po*�u���UO����4�j��-��ux�ţ/4�H(���s�U62i�Y�OG�E �QEu��Lν]#�]��J"O�A
��f�Q{��&�D��da������� $=��'�G %�|�7	�����{U�t��8�)�6��'�
�)�{�â��?6�V���Ls�%�89|T�Ѭ˔�T��F�	#��r�;���:ɟ,6���8T������u��3z�9Ņ3XP�%r82xg]�^���V	Q��oa�<Ly�ˏ�[��6�Wׇ�>3����K�]��[�����S�!�����8J��
x� z��m��<_گ�+�}�9�<�ӻ�q�"/�g��F�%7 ��7��%�����/r�B<��;+�w�l+˾�;���2!�&�Sn1[ �1`c�wH���&d���Z
�F�Lc�2v�_����K�v�N`�֯ԩe��\*���=���Ͼ��ӟ_[����6Mk��S�	W]�����>��{��䶱������3O����4٧,��G�6P�w6(:���ՁP4M�=.2$O���k�h+�r��h���Gj�����!����tp!� ��l�%�i��V�w tN�u]fJ��r������6����s��[�h�/x�YH��n������S6==��/�&ʑ�[G^Qk��O���.� `��Q"	�=ͮ�%a��a����u��3�R$g�ۃ��1 =�`Y�Њ4��<�v�m nEND�o�qΎj$�kw��}7)l�W~�פ����,��@g���8�͉j�H�;nc���ӰQ��ep����x1�L�/�6�����็�nj֐�"��&&���>�������P�ZC+�Pw���F�!����	>Q�p��M�vUni��X"_F�����]�;ͣ��/���g>��tk��p|�qTN�o��s%�� �~���h�l�]����a���t �}��;U�����~��ܵ�?������c�Bi�?J:���)k�b�5nm���޴ߤ���^X)Ӹ@/���2n>X61]��#;hI"B�I��o[42LC[�9e�R���L"y}�,�)b��c!��ݴH=��׉����uo��/>��똜��v{�3Si�<�y��Ɵ���Lp���˯�ZB#����
*i�.^,���g�{��S�;IJ������i���.�q� $�N�w<�5��N>�VD�����ʘ�V�`N3�����,ٝ_�7s�%�t����	�a�&ux� `:����$�G_U;L����f�� �����Z��SK���ī$Q�'_���Fj��+gĦ*��9��H̛��~+�8�uZݷ��|5�,�bg�Ƃ%�◶�#�i~Ni�O^�<HW���]�k����\��VE+�����FB�����*�Ҽ���s7 �-C!F� V�։���ǿ*(��֢�P�Z��U�P�/���D�&�w�+��g���O�v��k%����%��x�E�
�@ίC�UdA�fs�2ոvt��f����6R��u�g�$f�3*��0�`z�n3\pO��者�˰�o�����y��޸9.V��`��Ze�50g+$<�^g�#?�5��P�0�)��@b�������F�g�ז����UF���R�"@S_�1��Q,�18�/�OA9�mTA�H�����"���1�0J� �zC������s�B�3ɬ���*��/[燬RD|� �Y��u�@��N��H7'e��T�����~�Ds{� �>��DW���p75�5>V�� 6��:ׂj�cN�
Y�C�����%9�3�ѩN���,��3j��fh
#@��@K�))	%C���-5	���0/�$V5�+J5�Z��Qk��HG/u#�&-)��!=���s��U�n9G���2�8�;:I�<q��l�
�sS�BE(�b`�6j
� [�$�e���O+E��6A���f�����s+��fe��O�쎹�Q�M�OP����B L�JV�xs��yi�w�;D&�4���j��,w��N��Ogm�����BS���\玛�f�<��H5���1T�a"��2r��ٗ�!h읇ve������B�p�����)5�^*Ϭ�����k�V.R���~O;�K�/d���u�Y�,��,_�;�M-�K���!W�C�Z�0~Ƿ�����0!�e��EûZ��nc��S�dD$AڀoܬP%Ǡ�*!�.-�n�]\G���4�e���0|��29MC�\aa�>���!��na)!R�V�[(��
1$��,C�|�:?�p+�zD����׻����gԓȍ��'�[�!(�iu5d'��x�;�`�7��*U �0����䇵BLv�c�B�~�R����CJ|?T}S�ÓP�{��Q����"x��}��i⳧D�Cں�/�1�#�p��[	�1Ty�\��G����֘XX ��g��z��i
���je2\h�dR�����RK2���+����	4g[K�U��8����Bt�[P�������ѩ��}9�w`wiw�1�L�#)w�u��1'�4�7n�1�[98�
����%fL�&& ��t�������[�K�%V7�:��1{�')z����mxiOlFl�����3�^���2^��
��Ӣ�7��wEHG�Uq�jO�^{�54`O��X�&�R�fTH�t��Q o>v�'Ĝ?�X�-�㇪��P�EN�����]
T�v��][��s��\���X�����)�4D�;�����㳯� Wim�'�5���Z��
��X���X�g��c�@&����@�= >2�,��QY���"����x�#d�5�q��6��s)�u�oO8�jS��ݫ�?�4z��Ö���D��Ȅ�+*�s�V�
�pNg+_%�o$`��Y'A�x�VY��J
�Q�Oꬒy�B����Z�@�u�N{M*7@,�Wd�s9*|�#~b��a���+���;H=�Hf�K!dO<�&1~�~�u;S��h��XL�;Z�c�S�5/���d����t ��oH�t���*5�z�Ք�Ll�$b�<Cɺ��񹈟ڂ�RT[��ٹe��ޣ9)dP�7־r龍��@���6�^~��%�ۣ�ҋ6�V�!���V���b��N�h�<� ��{�40Q���K <(��>ۍp��V!���𧱞ãOsE}T�C����)%�iN����yf	^�)	N�\��D������S�YQ?\�I�|�:��X��
έ��f]%}������JG�ײ�v3���s���p)�*�*ⱖ���%W�p�;M���j�7P.T�ٓ*1c�Qzr`�*5��Y�p��+��F�G��Øl���XM`�t�e�g��w�!d�������B?��� &������X �8��:��Ù�J8�/������Jy��J�4�9|�ԩVƊ��hT%��Z�kB���]`zi�Y�%pR�پ��l"Sj�̐��CЛ<�������Υ穽��uzP'|TIGD�\Aa��:[B
�
h���&݄���ozU;��W>E��}��-3p�"#$ �H�o�1�v�ł��^�����";���[2�:WT]4v���Q������ܖ2��QZy�L���~ez�R>%,O��c��4� ݧ�~��Y��M�S �O��髒}
==��|����� �M�f�����t$BÈ�r�����S��Ь�&�\#}�*%�ƽ�D5_����c�$�&�����t��t�zi�L��.��i����Qw�7�n�к��AVz�H���s~S��}��`�rC�9v��7����0u��<0uÕk��m�_'�W2��w
��T
D�_��2����-a�F ���{1>M�Vx��v�-����Qg̨���!�����6�7a�~�@`��V_�UI�����s53L#���8���0����r��d4o�]Ԧ�3g}�$\?��F*/n]��PMzzE�R��h���������q3�s(2yX ��-��Y}G��|�oJ潪�U�^'��0���y!��ڝ�;��N(���O�3	�Ѱ%��|8O�Z���p�z��֥#KQ�Q�qx&|\��h��˓R���GPZ�-?�ouXX�����4������"���n[oG�b�W$u����/A�ۤ���3�fFRxK\fX'u���O�7�����Bp϶k����s�Om�	���{|��ya9�jN@�,
]8e�?��3��nxN�g#��d ���Q�Ϻ2���&,�*�B�w6�QsE�&�-�-cI�����Ǻ�g�-�8v�z�ẋu�b){�bm�����':�Ke��,���Lo�7���i�X>r�G5��s,�kʲ���_��Ȋ���I\�p�G~�4�2���/��x��[�@�c����1��-�L1�� Ղyu���5��1�����6�緍?���SՐ��͐�v9��_y��7�έN��*�:g\�Zt[�?e�]:��Y��XD;%s�Z��~�(+���o�rp��v@��� >IثqXn��CC��{����Z���]J��<���9$����nf]�h�$���hr�r.^��m�k�2�3�&�T�K�P�kk�C������j/c�f!#�@�!{���b(�W�p�1����/��U�9�utn��ek��7��TH���0�y�Ob{��˧"�м�qA^�>��g���p�W!����PS��)x�KzuB��sO/��^Ur�TͯS"_��!BH�>*�{N����ܷY]$�&�W���p�����sUi�=&� h��K4�/a��>ߩW��;�56豺{�&��������H3qh��1 H�������!LA�k���&��)ٶ�UO��P���]m�&�����Su.�+U�V�=H4O���LJ��-K��Cz�̙(T��E��&-��ծ��$�����9'w�_I?�,"��ӌB��a�N���)�5MWr�Αße�Q���W3��X~�HB���k����������Z)����m�Z6�j�#)�������2Hl��6��� �)PI�B)	5J4��G�qZ�;�q>�fe��Ӂkr��/�%P�;�9"ZㆲwV�r��|�ck��C������'�
^�榽�(�L�>|��+[����˄Y�D��s��q
�0�Aߴ$��Zj�A�piJߋ�ĸ�����/����^ �\�;�{��=�ǒvs�.u��m΁+��+^
��c��|Y�H��Pш�";s�U�b�a�5Y���g��T���i�v@j������5���Ϣ�-��yE/��w�N[��b�g|��G�m��p�
.���io�C��"`���� %�_)�#+�;h��ׄ����zk��Nj�g�e�n��F���xe�D4���y�	J�;P{x��{3��";+W��˦	0�9Z"1j]��C���$x��vA��`���Zh��kh��-����Dl�ޭ7✡��xJNwh���V����̈́��5��bɦ�A͵�Qtl���	崛�K��c䲕彷ڶ�Af=��~�}�t�K�y+�Lg��;C�	j����k��j��Y6�^|�����mZl/�6��]��ҍ�]���d��k<���R#$v�K�yiZ�J|�\e��U��wz���mӐR��ʎ��/�aG
׈�P�F�(��3靶pC0�����;��,ʓ��p^�Kt
��r҅<�Ye����W��$�s��H������8��d�?Z$�� U��L����U� 7�#q�_�G�}nʢ��-�7;��-��Y�68u��`��Y�������ݒ[���LE5#aD��t���)�h�*����*�'�NVc4���{Z��� �Hm��o?]H�8>7��C����7�vq��N#�9(��'m����8?�iuK��=13���	 �}�KϹ���}�$��_�ԸU�-P�S�c��� �g@�p�=�G/u�)5��?X��-�%��r~?AH���0��C�Rņxq:�p���}6*b%�z
�iv��^$�,v�$��q:vU�����kB	�$O�<gv�O�]�M�c5����g�' ��D�#Ф'VC��:�n�+�Z`)��Kf1m3fS����3R ݍ��opGg�S�9G(=�{�?��A9([����9�í�R~���j���ߵ�����ø�s	�֖���&c�ɆTB��8�S��e�����ː��*�3�Jr��(Cq_��SMR%K�˝A�jG�u�"N�t$��x.4�Df]?�-��{ Ƽ_0�E}p�������s�NL$�U���y/�=Uy6oIĳ���O�;M�QVp��!4ř�@��y�燧��̦m�������"�Z2aEhc�S�8�Ѐ�����iA���ȃ"BO��*�G$y&O�9��D'M0�r�=��(zZ��ǜ��0��o���+��w�l�l7�E��,���N��i����ʾ�|�-UA�K��P��K�z���j�o*����՗��U�o��wz8 )���X���w���1ڌj IL�i=r��J1%Q���B�����"zI꣤y�yo�
eΟ�z�">����$��h�Ѝ���%g.Vn#���K�N,���b��v�*�f�W7!��S�e2��jW»Bt����2{4�\�
�x�����a�[׿��AMsЀ[��<!U���T�� 1�,Y!#J%!���B��7k2��w��������u#V�l�o?`)d�<��[�Yg�e@�_iI	�e$?EA��u��&h#m�H�v`¦���d����ܤj�j�
�x{��|:!ι�G�D�P+��+%.o8a�T�Y��S]�e��d���������K��u|kh����?��d-����{w���'��lwM�F-�L� �(&4(;��n��5�bx����Y��&�8*ǡ��W_Xy*+���#7	�u
Dq��K�|��T����|0���1dv�I͡�+���A�>��t�0�n������A�����|ٞ�$�R编�3&}��	Ł1ζ���x�G������ *y�l��gbY���0$J��7{`dØ�9D)|y��C9&�Q��Hu,1n�P��R��)���~��,i�"�A�y#'�
��-1t�m
�ȩ�nV�h�,�c�y.��f{q::�9	�.՞��E�9��I����-I����L�tt��SP<+�5�V(&�?5<cv��O�[s�
� ^7q+`4��E�`	����,����o�����B�X+����E���_�>��@ wN6� O�|8�y�d����͗��K��{�7�l�p�c=sn)6?vF�}qތ�Vz��Ơ��IT�&Bt�2�q��ư������"WY��u�!7��G���B�JD�	"[�c�rN�Ma�+\�FlY�f�D�|�ukr$O��<���}����	���N��Ec�8݁� u8�?4�O�3	ƴ�=��ތ,hv
[�7������N'�p�3���'���)h%���/���u�jH1p�j���6�����q@Te�5�M�P!H�O�ݧ�≔d�	�=ajp���񝂛��h�����)��+e���>C�J���x�Dq'栨����t�ܺ'�vv��Rg��h
��ͫÌS�'��MX<�^��â��)�D�
bͅ �ˁ-���N����~pl�]���8ξ*K�3�f'��� i��+�x,?���h	/n���C�_>�X�J䄿!!�!���1&��3�,d<1F��]*Z�Q�]���CY�:�}��A��F������x�_�"����}{�+V��	�?Հ��װ-e�%^ �ϋd�˲G��r>@��c[�,Wb�cO�L؊��ٓ����*�a�W�Ft%tt
���RP�yi냷�4��\���Ĩ)��鴧\��w�朇���)�� \a��o;�<�����&9ؠFʂH<�n�����]�/7��T$5�ES�n�{ ��;8dC�|�Cfw�d��C� ��s���pz~�����ߖ,d���7��T��h�C}�r��L~��$�&u�38�� ��9��-D;#S�v������54�3��A���"�0|�%~Y�2t�RIS�cMo��!m��4	�´�v|���?�ͼrH{�=��G��i��w��N��z��w^w�����@a6���k1�6M�>T`�����8�u;�7BF�;Gs��-1R,R
������y73Z�]f������0Q����c��D���#QX,����Ya���i��Z�k��(C�[�9W�G5��- -�SB)~�p��N�뙷�����ӎ�o`����wl�$x�����g�Zr/� :R�
���E�Y9D�ٙ�AA=�Fz-��FP9����x�3o��l	�a�f[:��jo
����R
k�ԟ�����n����gp�vn��a,~��T*G�S�\�<]��'"_6��bST�0�Ȗ���eD�e��ާ]�F��!;�n��~Q<Ok(V���n��4����y���M`�n�x��D�����љP��Yo��+��3�+�|�U>�'F���/M&CM�`���8��I�"3ּ�<�*, _dr�&��{����+���J�A�
�!��Gjukؓ�	/���ۺ+�|.s�@�>ˤ�ܨ��t6J�j�I7VO���E���K՜᭨�]�s�qT�e0!7�o����	6�<�u�	�y��OL��(�k���%W=�(�����'�{��������Ĩ�5�F��dwp֔��
/~�b����kWxU����$��fNT�q�3x9;���XV3_������I!I�ftEHv�/�N÷�QwT�̖��8'�^N���D���,��>�J>�]*�E5�J�r�d��jG�y�zh�I�Ӝ
	�t|+<���Ѩ�����0M(�Ya���{�tL+��poOפ����/�l�����	Yj��O޼7�9Ѝ��5����J鄶�`[�Ǔ�Aq�=Y�ց�׷I�A�*�ܯ����gG*�;�Ex���IN_�:r&�a�z����.�9"/l�"�?yE/}��K�Pb0��z�!i�\�YЙLԨC��%oź�)r�5��3�p%��>xg6X\����M�zF�
 �ҁج*G�OY��W�P֨�è��MCt��	���S�ɘ��v��{P�Q�nf:2��Y���mGIW�&\�]��A;oaV�������0��vbxB�=u>?�+M��f�*�<Q ���-+���0�g�{�Mx�,����'��P��$�.���W�i�� \	���SH���C?����[�;>(�`r̠C���%x�u���N�_�H4E�3��.�����'�VT"P��/U�Uy�1���B���!�eYɅ�I� 5n=/xC��4 _��ʞ��oD,���@�6D��w���ì�dC��n_��us���X����®)���uy`��w0�~u(��˱�����Qn ߹����b>�s@.(�ih#���|v��>��A�`Q����ō�JO��Ѱ&`����#pY�fŲ�K�c�b49Z�m	C��͉���-�T��ϧ�I}���!M��KcѺ�Ѯ�� �"A���cs�̮KLELAKR㟜�Π�M'V���4k	(d1��ѭ�k��#���5U��'����*��|4�w�q|�05�nV�t�>�����Z�������)M��E�;m�=�&׿�^�N41�I	�,�#���.��71�� !�<���C!"3��&��~��hǪ��"��m���tN�4�L?�#����}�ң���n�����M�8<9lIk?��V�nH��݇��ꂇ��v�a����A��"��#j���5YW%h�/NU��pĪK9��D��`���d�^/��,�|�A4-���=��+�LL|�ݟ��_��2�?�K�{��\	����SzlH�u���)9R���(�v��7Y�h{w�9�P�B�������
�Ŧ�eG��\��L�p
�/���w	,����qNu~?KW^�N�
��
��I��ܢ�bo�3��!S=EJ��f:HxXV8ظD�$���.�W{N�E�s�ZUc8iI;��� [�jZs��D~7J���LeNZ����n�u�:�mP�#����(�f�B�_�|TXҬ{�W1���K3�4�\�g����/�ˤ��ϛ�����I�KeU���ȷ햐(3�MF_It��Z��[���2��D������Yx��-t������#�P�j*@��>��}2L����όmk���!�΂�$��>�AR\ι���s�l|Ƿ6��0�>��Uɜ0L�Z�֝��T��YS��W<|<m����7���/�B%+Q	Sx�꙽�$^��ԔX�,��&�E|8E�H��{LORA����Rc�A\M
;��X�3��W�K/��I����Q�t�@�����>��^wQ/��n@����sX�ъ�s+�����Ai8�J�2��i���p�Ҟ��VRa��D\�L���Q��ӾC6K�_�}�4���'|�ɑ�x��^=�~O%��P+���z�p��s�����׸�k��K���h(�����)��)T��0S��S��}p`E�xu'����Y�:/ߥj�~H���H�#0���o��*	���6ac���n��Q_�� ,/�}N�q$���zʾ�a��~���!-0&pn�(�aÔ���5����i)z�\�@��#����Q�Y3kC�ի2��R�_����m�1��v�K�̓�?�7�\�&Z���85t�Et?^��Ez��Ȑ�bD9�iu��@��OGu�Hˮ�Yx?g{g��I�q�/}Z,Z�|�zl����ؽ�Q�a��
��^d���>�'�����s�t�H�����g3�y��#s]��h!:z��2��"��4�{�H�;}M4;����K����K����$F=�(�?�/��}W%�"��om$ʽ3�TLi�D�{�z�0^};39�\![陞t���I	�o�;'��+�Ч4�����)�$gز��k����A	9�BQǈL?��t;q�r�`�g����	C8�'WK����Q����%�CV��o_�'���-��;UZz�P�O�l�|��ʢ߄�
�}����I*�t�~���pG�lT|%�	�By�F���6<��8��	T�zQ;+x[0P5��梢���L[�܃%,���(,u,�	>�jU�G�&��Wo3�����}�r#-a�>X���A�0��3�|�狊�FQv�߱�����퍍����{�fz�!�}��A�K�z|{�?�~�(]�t7��e�+z�T��AR��E���I���/q����_��b�!����ja��|֢���A�MJ����Fk�E�$# �mRc����),k�D�m1�i��3�� Z�ރa؜��v�J�Q�L�Iƛ�ә�Z(�ӍU���\���8p�����RӘ>L#���Ȇ虵h �Ŏ�T�����;3`s��@�����v��E������6R ���
6�5`�H�%ӓw���b�S��a� Ԃ�k<�c�^2oD�B�w��Ӵ�}�"r��q�Kt?8g̎Ր����7�N�~�3$�U˾"�:��}�3U��>�*�h��)��.ߏ�y����)�5 �-_�4P$�3�2R�R�=��?RK��.��}��yd%�i������c�q�?~���>)�y�,)���K�Ypb �"ʦ�Ki n��ӼGC��Hz�Є#����b=QD���M$~6�<1��F6#-@�U�-���hg
H���Q�ܴqhq��h%�dZ��y��t.��A;5��6���D���%s�SC�xH�'�@VI$�K��׵��H�z�Jr۾+�*�)���.���m"��;G ��NMD����q��Gp�( �}E��A�2R�34�(�^T���,�)�vSz�G�*��|,�-=�g�T�� ���w���9D�Zqy����ЋzYH��Rh�Q��l��;P��*|�|�i�ڻa��g�kre��ycU�& 9�z���}+��>C�:g�<���e"��e{kL1Bݼid8�V�M���.�v`��j�)A����P�u�����c�Ь Y�S���9����L����ԉ��S\�;��E�ÖAQ���1!��v#��s�Dx���|�=��üp������g�6�D�T�
��W1����.�M�������Ed�w�c.7���r�P6�T'D�Q���b/#M�s�>V=k�DUzQ�XWaf����D����0�A�z�R�~�,�{��І3�!�k|�e
�ݺ(���l!��/�B��!G�#1�z^�S6<��������5-��XM�aGʚ|�����AϘ��S�<�W���lں�XvV`T�jvj��`�D&�r}�����>�����q�s��/�~���p'>��R�M?#R�
vJ�	�v� ��WwJ���v�.��4���(�]���T#���[�\f� mM���J��Q.�h��'b	����8�YǦq�;?�̕��s5p�4�"���P��1����Jo�D�ٴl�ny�kL��Ųdw��x�rw=՟�>�u��p�?���& !N��P=MFyP{�'[]�TKs�I;}V���c%�[r�޼y���z���%s@���A��p��!�)嫃c~���M*q�f{mMnwb�b���~��l�A��[�bHܓ��
v5������"5	�����Ѓ'���J(���$�q��gl�C+�����汣�(X*c�o늋^�x8MCg���5À#�bj7�"�<�|��tg`��*�����jam�eb�*.�	��#�"n���gv�۹rq٪|�Dn���kizѲ�o�Z��9N&7��*C��P��<P��T:'��"m?7>�vz� ��;��8�t���T��:j�F~ kj�Vb�ѽ�����-?(�둖�L1P(̌c�^|k��7�뇰) p""��ˌ'f���Ot[�(5�4l�C����)H�6���}�~S�-c/����$��X1sȨ���E�]�Y�Z?DqY����R�fY1`�B�A@"g;��F��+u�|g57�V[��)5�q�ȁ�7�s��s�6�r��7��Y���Lr����&���8���ۑ�ɕ��Z�M ���jb$pCj�m�E���������L]�#���x�������� �,����Ӏz��Ղ��*���[�98�q��8cJ��PE%$Lצ���u�ȉxPw�o�k��'����-�b@�����*��:&�M�?ǿ�Ob1G�����5����i�����)_�ٔ�?�!:��O���G�)s7��Jf�~�C�	��ؖ+z�ӣg�u���hj��h�!}Kr\���]�9��wn˜�k�.�n�A0Y��k�Y~�tX��@%��!H���R�J|&;�F��a
C���	�\uG��x�m�3�W�=����f�x'/����W�|���0e�o��������c��L�n�<ϧ�����s~�7	b�� �W
n+�)�D!3����}t�I��?�F �Q�GDW�[
�(?c%͑�jc�b���y�  �C	�� &mqv�%�R�"Z��V�^�r�HO��Q]��"$�Ʉ2��H�G���5k� ��r:��_�|� ��,����(M��m(�Ib18{0�1|3��f�j��Cqq]�f�aG<g|K��`��+6F�N���PI�a��������]<*%z��U�F �!*�$hs�S7-�����[S�_�c��~��~�<({�0�'�GH�kH�{.�� xUAxC��OJwdD~���e�e�;['\
v����������0�v���i�z��nH�=U֖㉍�%ߔ���/���ka����_V���e�KT�ũ$�
A��p����s=��u�hujb��J�Y^(C����<��a��j��f�QM����'���2K�<���͘׎�JZ��f��:o�N����!��"`A0�X�����%�X��>���]-g��T}���U'�����>�� s��9�8�=&b��q�F�OZrK��vi���b�`�dW��Z�*bQ�׭�۟F{cj�W�)L����4s��~n�r��h�~s��s�O�+�5T�?������XS�ڱ��+��`�|ܺu����ߞ>Ru�����4�I3�"!�Â@�#��(�)e9C.n�M��c��bQCa6�ɆwP�T>�x>G,C��a�8��Z k?�o�V{��u�5�4�N�^J���(Oc0xص8�o�(���Ǝ��k�&�v��}p�� ��a!�������ģ3 ��b�tTJ䧥��EqB�����
,Y���f�5U����Ǵڶ��<P���jB~%R���LN� U�v�O ��đ������4Ϫ����JeNw�� W��Q8+���v n���Be���,u7��צC�|�+�Wą����'*׺�ؠ��>�}g��_�+}��$�*r�93�ę�}[��w��;�����h8z��Ȫ˜�1��_c�Լ[��; B�(D�L���:�U�@��W��#{�U�P�r���%l�0�������X��0��>]`��b� �V��4�ɑ��X�s=E'�(��������{���%���N�9��k�[�K��/��i�P�w&,��3��\��*��iR��-M��A�o[x`/z����s��<�W�������<��߈76���~>�J7a�����VM�=쓾;���/i�b|��4X�5�uj8�y���]Ý��bCj-��v��.��1��Z�`;M����-��Ť��J�`��'�5��v��l��<˛��F=��lg��@Jϱ@n��_L�1�u�K")�L5;~�Qa�N���`C�^�Yv]݉�[�	��j$%>V���2�K������ń�H ���"�{��zL�y��$�ebH��C3�8�zö����#x)�!W�b4���|O����r`0�Q�s�k������w�I�t��y>M&����Y������)�� �:����/�Xƾ��� �d����d\h��'P1��[��p� ��)�l��\|$a�q\�=�8��^w�����d����{U�a ��4��5�2��㷟)������)*�;������a�#R+���?JyZȯT���
�2��B�RR��%Ǐ�(QP���D�0��3R֯+C+^֗�t2�Ps�p�3Q���OR��=�H	��G��IW�--��>{���e����@6�h��q�d�i]6Xl��żn����u��u�Q=2�@ZΌ���~fg����LAQHpYs�w�W���"H��EH��
�h����3�U�[�+�F����OH�&�5��� �1��9M�y2���ʮ[�i�za�r&g��Q�_�E��10vD{O?��������f��!zp<X��V��>v�T��kܠ��'~�V=�d�^�%��eT���ӂ�����+*��n�K"�p7�蕡��M�Uo���2�� (=Yw����W��@g��F�F7�TbZ"�Zx^˔���]'_����x���ʆ#j��Z�~�@�u�\g��$m�h��@�9�f��v�����۹_	����0r(l�(Ϡ�rW��X�;�.�}�A�Xs�}�w�OF��O��o��Vuڧ��ŏ����m��?>}J�������є����m�%�[���� ��m�:��ꇉs��J�P0˔o�d�p��;F��<�� ?���y����sk"���b������;�M�\~���&�9�m��;����4���~Y�N���?�ɐ;54��j_;V�(+�{��4��x�nm$��/���S���c��k�g���4�̎os�gǽ#�2;@R:�  ɖć�{� �A���0#���w�tBxL���[Pr�͍+0:-�Z��Ah�q��"[!�t�F��(,�]�X@&����L��i�ֺזY����SHWf�^g��śoU��7uƛ&A�]Ң��K��IZ#f�2x,�mv�f�.Z﨡��Y��~{Ox�&q�&�	�7&0Q�b���C܂�Ķ�Ř��b��24-W�ק�hY�C�YXέ˜�V1w#Ϭ�Ɠj��e'f��4Y��� ��S���?��gV�Μ
��6�vr������⊦2 �� 4���7�� ã��O<�D�Z1��M"�24�V��Ns�/E���������|7gH���2m�Mnw�"3(�_���2RT��7N0��/��jIFވ��A�b��BZ��k��[̣X�Y&Y����G�b{9������o�7���[��4{Q���t���C�L��C�m�*5�9����p�����h�M�#�Q�˭����{��(�<Y}��b�]���rXd}����x6�&��ą��D�ۄ[��{\�Vw�+�8������IWT�|��ߒ����ɁV�]Ű4H~�mN��]�Ve�a*�làO킢2�n<���$���� �Zr �o�!tsc�R��tP�������l�L�@��]?(����C�,\��Qo�ɯ������ V8�Jk'{&����uG�	J~/H�y���t����y�_|���׆�}o�g�#�*"������Co;b�+zJ�%��֢�a�f��#6z�;B��4�|p'��~:� B4>4����L%BYM�)a�?����gB&lbNR�*�'��)�&��W@�G��%fZ0��,X�YV�ypP���1µw�7���9�,�7�	K�P�!�+�⡅�m^O�*
n�	�s͞�w4�:3��Vqvq�ռ)��0b
�A��� �}��,�/ �ה��-/F��#�Q[��E\j��%	W�w4TJqͱV�"ڦ��ºUW�v�����S��&��U5�gh'�u���#�_�(��1�;�����뎫6������Ǳ��� ��<ʥ�����2yF��E-"ߗ���+f�}���k��P�����qH�s	L�c��jEy@��JN�."e��}��n�d�tnq�g�>�����T����K*�^�[G�<��0�bo8�uP�,���U i:^D/T��	 �t�5��6�Ы��xU}�n\f�@{�E�p��޹l��%F�DP���7�'��vV1	}=q��j��k2��"�(�_���r����P� K׫aL��j�|��C·����N[Wú\��������$�{Q�0;�-���_k�05���`�l�W�kD���Q�'�����O��e�7�4�'��Vu{�S�����L�Q�{xt{�d�)=�LGo�X&Q%6��t�СJ"wi� �e��l���i��Dy����h9��S�fl��Y�L��Ϙ�Q�#w�(����::��D�H.c�+�.j�+��Gؓq
�"���c���"A�4�#~@ǀ:S�2�F�6�껕1[�D#Y�)I�z����M�����.|:�c�lU4��k�5_V�C��0Uj%
�VaF��N<�@��PH��<��h��@pw���\��D� �&�N\�]�,�nIR���I������E��Y2�pe�e���R���sRMORc)U�]%)�FZ�Y�{�_��M�_Ï
H��%s��k�����k�P���R�Z������s��hL�U�ۺ�=*@�RQ�VX�I���<�+u�7iK�8���w�4,��[\���e͠h�~�h����y�}�b[cUB=�㎝u�a��Y�:.����.s�!��SZ����!*U�E<��q~�L�3!������i��k��0 �=FA%�Ɓ���f��C�v���!U����(}���<p����h�G,1̳���4$�Y�y���U�?Π%~�!��(�F#n���/���x����M��.�0��x:���@�}�\b7Q࿽zƟ�Q�svsg5E6��８p�<uU,�Y6�#9�K�M��L,1\�O'{�f�]%��j�c���Z9��k����@����6��V�"Y���;�_����i E �ؽ:5'�	hV�B6��El�Q��	�$�-��{����1u �C��uER�}æ:W��L!`�f*����5���p��"+����o�꼃dE.�$$�W{z�>��-��-L���e���������l_L�|��
�'�����1���5UU��nq�B?C\H�����ށ�/]�(�3o�NÚK���n�p�=&,e��b�ǆ�BDu�ߧ��h��|��쥿��#\�S�]��w�-F{�+�v\�#d�I��ٳ�hhq�ƤO�?��Ӕ�i|��~A���<��L�6Tl��ѬB �p��t:h��M�4�:���h�E����d���o�87��HQ	�PR(�N�����B�'���ظ���@�E��Ϣ�?���Ho��GU$�Np�ۼ���_|�#vے���#�=��Ψ�?w������`[�p �Oi�g~�hwJ��wj�?����!5ç�EZ%Q�G��|G����]h�ѻ|v�7?$�$��}�CX��"}�|㊑������s\/*V�t��?Z�E�^)s��P���h�R�r�,���{�W�7CS?��b N��AP�l.S���'s�A���UL/Oy��4
IWT}��FF2\#����Q�8�/�[ˋT����Js��s@|[����VX�7�{q�U���뎧f�m��VZ����Gvh0�]�\�&��J�]W��n0�dL���#[��5���j�j�=P?kc%�ы��K��z퀰Q���SIk=�4�C������%U3��/�����Է��'w���&�`n�2vv�@Z7���I���9֛�uV��>��
�E��L� #ؠ�(�O��g��I	��\���/!�5�q��4C�kKcwA�Cnt�K��N��U�k[�`H»F��!هU�{���LȘy��Gh�Q����3V�g����AwƍU��X9�z���l��o��"@� ��"\�*��k@����8����Ny6��˯�msd�  ���S�]�L�Lh�
yͭ�tb�MV;�^�G2��ξi�B���F�~�_��(��,�ho֖s�����]�a�n8�Թ�p�F(MC��^�W��Y+|��E�E4]�R�2�N�lv��[�S�]X���bC�h;KVF�y�E��_�
-���☄q��n�+�,�9��C���E�P߈%#���m`��vY�Y~_{�����	����]>/	g�㾫��?4�F�cA��IcPwh꿤1���as��Db�jA4Hߣ�C��I|���}?u�	/z�"����n�W�ì���B�$.������Kbԕc0t�6�F"����e��P@�L�[u88�q1Z���7FҸ��Wf�!�^'TؿD�8�'� ?�0d�$�3��\������'	Jz���A�:P�@����B�z���_�gȟU?�J v��f�W���o<n	s�J���R�3�L�y�(��F��GIҜb�����Ú�LwT�w��^[3I����[�d~DS�f�s(z�@��&a8�kV(` �ϣL4���H�|���$`��ռ��%&O�|?L	�G�u%�z��r;)8�-�@����=m_~�!���&]kb"+[_v,廩����ʚ��*~7�����7Kج�Ć��f���)���;2��jl����$����R���Y��)�c��6�ո������Y_߆��&|T&M`��˃�K���ܑ�����(���E@;I$NDYK��	�Ce�{����y�ȃ]��py8o����M��c��L�;��v3@���)̏*C?	َN�h��?r�\��DƶS`��u�������K�e��178.Y�Ǧ�^G�hh����bEg�1Z���D�����&��y*%'O9%�m�
T����3�4��k��5~�^�n��S"������X��C`D�, r�k���E�C@@�Y�{�L��^��L�G��'�
����_��G�เɼ�&��O��ꫬ�B>F�nw�}����ф�s)�M�;�A[6F〇�dx��J�WeN��N0X�y��C�Xw-���p���K!����� &�,�i-E�z����"��|���6���*���ҵC�#����cj�z1�UDv:�8�k�jԠ�FI0��v��mǿY����F�)8'ΐǼ���o�0O%���d{���ɋY��6��1Gxa~iwԋe���\�r/�i��l���к�	0���v���R48M@뾽0f�
�%�	�֧_�+Sw,e��`Мu3wN�j�#R,9�,d|�����v��L
hU��4���ԛ�r���'�S�	B�Z��i�2��=�ӧ��o��@�	G�>�s>ۆ��G�6����G���� ��6�tsx�\�X�l�Y���@�OЁF�ph���GK�{���
]Jq/�W�R�:4�U�:��)�߯�����)���P~j���:�n�nनI&��U:ء���M�C���kٹ���o�z��:�K�z�sr��|R�F �����{ţT��ש�ra I�v�#r�\ؙwk?A8Ucg��-�������D܊���A����=~��2�54|�{���q-��p`������p��N��^t��|*v��H$�{�]��½�bnS*�i�=��ڲ�¿����|�y�N�@�g��/y��}�ɊD	��R��޼\��L�C9����~~�q�d��-C}uHI�U<v�P��|�v3����U���'��fh|���E��&����:�nK#��=���`�J$g0�s��|SF~�:V�X=GR�7fd.!�ܶ���H>3.rr̕���k����Z�?N$�v�C^RԊ�GnU�a�e ���ϥ��}����h�Z5M�L��������I"Y��������7;��y�$��s�L=�.�f!>X�U�@(�C���w�}�RyĜv�wA�?t[^`��bb�jA��v���Awv���4����Ѧ�6f�p�f#�A�[���2\�T7E.��Ȋ���P�~q;�]�Ư�rx��,n4fc}�����=I� +�FiYh7�<E���'�0��9�j�Fˡ�C$zA�ź����o�(����Z8����9��l��)��Y{vJ
c;�(,��_F2GOq�EHQ��������t����O�����b�}y�(�$��e�����*��,e�{��4*�k~��|6�V��V�����3py�\�q�C��<����@�l�c�6��|A�QV��l�)��ڷ&B��U|��[C��X�}�b�@�����:֢��7��b�Hy�YB=�S��N6~���Y�҉+�	��A@��W��h�i|C�|'��#�ᔣ��!S��	6��s����F4�.�HR��J��� �b�Ad	��)�5����`��-u�Z�e?\���_a)�v}��d���D-\S5?2T'� ��;�0?��v�&� a��o�@�1w�I��2� e�ccT�T<i�`0������� |ue#VTU�e�q��܀�8Y����]t����!,NF�Y=j��̍/�[�/��h��5������LB�֐�z�i�q�$��� Kť�3& ��c�unC�k`\P��F'VO#8�K�B��V|�]clαhjʩ*��X�+�:̛�3mF��z��y���a��~�=	�G��dɺ���)������W��bE7�:�E����������Ǜ�.쿠�R8����h��m�խ�m�%�1����1,��G"�J�Pߠǉ�k��@#�4,bYo4��fͥB���z�j/�Kb!��5���{�v�O���C�,V�M3A�0����5#^C�t�`����ho�z�D���9�x��~��&�)퇪b�X��*_�>��iq+�E�t� l�V$���ٵS���ï�F�|���}�0�9k�1!z=�̜nx/ �o�' ��탠���s�%j׎WU��8�+�s(#/�� %��1)�a.�h�)7 ̔ԃ��g��_��dU��K�&;�wxV�$l*�u���4L�^���-c��H�(y�^`<�R�h{�w�%Q�
�2����	`�J��fx�+~�_>���E��78�@��\�4aD[�!����+�~7 j5Ѓ-�Z�R\9�Urf֤c}��9�T�ٴFl���W4�_�Q��6,(�GA��MM4�],��}^��k�^�Yn'Xh�s	�c49��i�Mֆ� �;5�s��{��hW�*̗D^�{�\�+�a�p����M�5�P�>v_K	��u
���8'k����xI�J���*��m���T'jA�L�[��f�=�t2��CSC���0^.*[���xë ���E=�� ʏf�P��ٹ5���J`�	_?^=��I�A�~�!���g�Z�nv���"��\����3��:|�f�$�/�DJ��-�"&VA��{E}I$o>t�m~�iSN�4j��	�G�g5�ū�g6�ns����g7��⼙�HgPy�$}6���ؾ��,��?~�і��8���b�T]�&�X����y'�g
�Z�H�;���1&�s��l��8H�`�R"�Vf��2|�5�����$�����y�8��䘭T�uK,6S�(��w�\�pWJ��q*l�x���١[��Jv(hi���y�k��3�%�m�2�"�]��^��	G�()3�8ao�*5�
�|�a(�d���(�̀VE�^�p::{W=/�ؗ}���j����a����5W{��x�p)�ZX�M�et�'�$�ǫˆ'8�%0I�&ǣw�׼��u���~˕��a�c���:�(�Fu�e�g9��~�Yt����b��xij��M�y~��>�Ei���~ ;��(�A��{�ĨJ�6;�pe����HJ��6,o���+�>���,���hGX[�^�m`�)-���2�D��AO8XM�^�:mH�
�K���-�>"��:3Gj�!]7��a.^�_�|3h��)VV�^���3��^.�����
�dQ�g;�}^���}.AJn�H�m�� ��9���TXs�3,S�X��Ǐ5�2��q^�:�4��V[I�!�a�ݝ�9Y 1a!�/ݲE6�Zח�0��IsO�[�1��Z&p��A[A+���_��v����)�
Wu=ꊓꭨ�B���%�]�BF	:a��q��^�5EW,��sy<�;xYv�
[��*�yl}Ml�:�Dz���K~�P�8pQ�ow�1_�gP ��h�΀ciOU�5���*���=���/f�����o�Z��΀���n����W�|�J�|��������M�����P�����zC^���
b3x����̝����7�|���>]��~Et��m�ٌ���!<9��"�U�C.m��ԝ��o�U��ޯ֥�/�6�oV��}�X���Bu'ڀt�T�K��󙩴 .`إ�6�X]�r�9Ί̰���\(�N�I:
����+�rv��J�z��a�H����:�=�W�"S1��-��O�j�~�8+5�s��(�Ұ��3	G��@���޺����j����p����[�v��*�.)_��X�۪q?���l�sU�Y�
O�u�I�����d�S�@�>��������Gm	ۘ��ʛI��֮�s�[�-s��qL�ݬ/4����b�ku��>�� � ��]�@R��:�r�
�})�p���0�Or;P:��_\�$?Z�L�!^��jk5/qŌ�~^�j��߲D9�_<f��QI�2�(��*+5��wA�
s����������#�9RW�Ql��mK�U,�+é���	��"��}���UP�L�z���5��+4,'�i7�=����MS�"�%��~�v�:�ړƼ?�:=n�34��i|&$ei'����j6�$�eԗ��}Tg��Μ������]����V�+,��Q=�:~9ߋ��}�ԉ;o�ց�;h�xYʘ_PGfR�/��owY٤12���j�[�T��<���U�n�-�ф��c:d�(,�j�8Z�Y�"w°[w��R�|����MV��m��r�&�ƫ�k~> ����ѱ��:����X�49n�t)��>��<v��4��$*حR�1��ˌv>\�}�ZGn��1��(��_vˌ\CQ�c!YwY$+�xë�ď̀��� (�f8�Z"��pqK�}r�d��N[�,X�2���02V�?����s�7�uİ��0��s�
��.�QX�hr�~����b}g����~S;�=���l�,=A�S����@��~#$ ��c�u_��}��ϞN�W ��d�����~yw?��k5���E�y�g�]�oyr�]b'�|�+�ʧ"����FBF�H�P�a#g1Wo*�!-�ы��2�sU`b|�����.�����{���Td���X�������r��ü:8��h�.T����,v�V^�I]@��Q<Mʆ�3J�fmZX�� �G,Cd�r����P~c(?c��(C��rV�W��m���ali����7�
����rr�iǴ��&tj�>���7���,}.=�%
�U�C���~��	�>R]��6���ߺ�n��eB($;p.��]Ͻ��+���߈�Z,�E��+]b�S��Z�cO�7=��!�~,?m�4@),��0���D=d�uN.!�����;g"˴/�A兵VT"�������n�D�܅"������y�&+df�F�*hZ�(���Ubͫ���M�l�Ts�HU�wE�r��Z�_�d[�ȋH$e��-XD�������\2S9v�2l��Ƌ?�H����K@�Ç�1$�U
|�qB/#�x�?{Y$8q,��x�?$�nq+�*��I�È(N�	�I� &G8�+��R{GS&]�-�{о/��K�b�_׌���H��T�œ�X}k�p����)��5����?��@Y
,eZLчEvt#�&
�ƣ'����EM#�~`��{$v�:^U65�MC&)����ET�s�������~ck��<�*7�
�t9\f�|���b���O8�#*�܉oA��*�v@�>E3�l~rk�	�q���|z��H\"��@y'��D��0!e^�������G³���Z+�K�a�@�3�W@�[԰ǭ`�8Uz�dE�j�j(��2m�M�ν��b� 4�/��.�!�| �誓�Y�m��PQ+�w�&ݕ�Xh�KqZ[��?\�X��k�:�9��(�=��*Mr��-0:��ϙ�=�ĚP�AՈ�� ���f��	a2�۸��~�jU�S�Pp��S��#���n�BML���_�rn�ʲ۴"����N4���i���a�ҡ�ܖTf�N������'��4���h'�q�r1�e��i{{HQC#����	�&h�Ec�X�Z^��In�r��z�o*4��:Pz�\�-L'�@��L�S��R&C-�����Ls\_ͱ�]�h��X���&rph�C^].��I�ll�rE�!J]�כ��Rzp@�S	�K]���/����ȥ�5�QW�7u��3}�q�U k?�
����V�>���^f��B��#����Mh�C��I�X����e8E�g��}X
��RÎyZqi������!X|�d�c�"�{c�3��9D�2
)�;(������HR���bȏ�K���m��7	��S 5����W��j�չ�\8T`�r����K��)Ć��+�����[f"ZJ�?����uffe�\���@�a���T��WU�M�Ks?�qu`NZ!���0�ʀC`�_�׋��K��*�d����x
ؚR�"~Kj�T��V���I�p�� Lْ}沎�U���FҚ0�+�T/�*�����g��������34���f�˒��}
�bN=om뮿�����C��a����Ǆe�z�$7R����!�	�tm6�J8M�]���̴��G(��3���ɑ$2����\�/zC�v�T8�d���^�(���9d��x$.��k�u!�����sL�tw��z����J%����%�*��r������f�賂`�M�k^.b��C@s��F=v��kD��6��b�^=]ن�u��y˗�z@m[[z�@�/%k���;��"~Tp�Y�����1���a����]����8n���j��~[0��(������J t<��M�3}`�\ɰ
�Ty�
��*�NԉR((EBm�3;S�^_,m��?�:D�4�L�}��JV��o�:�4B�)H<���������F�	�������L.�3J�+�vY:��T]ʡ��m^M��؈�f�Z�3Y/��6�{�3q��'�&^��S�X=��٨kYi,���xɓv	�Vj/<!-;�@���Е*�C���Xa���C�����/�-m(�ه�5K�Ì���T�t������x�1�xO�����w����r�_b ���-NG|��Tq�`�c�{�4�.���؄/~��J����_����ƚv3��l����R5��٨4��D��կ�r�7�# ��*���徖�
��-в�NZ��a����Ym��L���ʬ'��᭪7n�xMs���LE)�G�|�XƠ����c�*�m���Ӄ,��j�8�sq%����VUM���!�aK��%�,e��tFb.^�xVJy߶�\윣��H�\�Z��`���.�/l�`��8 �7���P�����r�ğ�n�^/�Qa��k����4{��֎m��:J��늼%�Ԋ����Ru�lQ�n���β�����/��M9^�����]�j�\���mY��h�D�'��k����D�(徴�9;��11\6�D�F�a\LBi*d�����g��f���}R��I�k)��"fV��}^ǻ]����ZA�P��pm�LmB���f��&G48O���N�u�ُ�t���w���H���L��\�k��N�X�-�����@凱,�)��<D�v+~�w�l�|��2�����LDӕ��l��mZ���'����/��齃@���C�Ǹ�57��=��*���6��r#��x0.��[����������<&:��)�a\fP�B �o=jF!C6���Xvn�!_}ٌ=k�LR�%�xAŏY�U �0��o�:����~�gXSH����hp^&1���W�C���t���S�-�����j�?����7rt@�\�p>"��Y��:��`׸�-��>��=ա�^q�����3���~fW��kr&A�5J���9o$��*oM������^g 4��z�������h� �&;BlцHě��6����Z��_6�BW�sj��4
f���k0/YԚ,_n2��d�)!M�n�V�p5n�_ �_��&��Ӛ7߳Fn�2���;x܅�d�	}(��'#@/�aO�r?ͅ�#����-t$m@]��;�!I���8��8)?��
_L�t��+1u�$ŝn�����^nfI鰃eosM]� $��P@����iA��I�S���?��5��O�B�(�\c�6�����ny�:�M�q�̊�%b?Ht%�Tܛ57��}��C�y��]�]�������$��QF��q���֚��צS���M����4H�E٘-��R�mIdS\��y�����ۗ��UsVi����"5��ZsV��q�a����ng��7_�������(�+s�/�ɐǭP G�'�U��i�)P��j�Ew��"���V(�g��z�#ٞs�d�x_W�GX���7V�T�֛��}�12fl��Ejc!�2}$�ӏ����ʹ��zjo�"{�A����A��g����k�RZ�ݠ�.L�S>�.�Yv�`��"�!� ���n���W=us��"�K�W�uj�Y'\���<���u.o��xx��r��(������S�|��<.Cȭ�V��ւZe��p���R�C�0���3�D�!؛ P�aC�u�?��鮎|y�0��@��y#�?��Ɋ�2A�����7L0����@*���0ܪH��R�{n����	�Wo��$t�3�^� k�2�NW�I�wS��YWw�/�,��\K������;>J��urJ���p�nK!=�G�cR	�?Q�fg��?�+��҃��O��2�\�͡%h:!�oc��3�Ө%w#�o�XF��@4�L�ڷ����6���d@�޻�-ўU|��'�i��B,0�h�/܌��1Ɉ�lPs�E�8�+��W�r�k�����ތtʩ�.�G��f:;�X|�
��2�乗��uN�~F5�i�wY��U�r�X���.���M�@��!�� ۄ~B|�������L`������\nw34�;������5���]Ⱥ�w�?�~��X/&Z �8��J�ZC�z�����ص,}I��m��'�9����S��T�
��z�p�����o�a��n��������$�4}��R�U3�W�P����b9FM56��'d	��>#7�뾿j�647;f��+J$�;Y���,��p�*�-�\Q��~z��Q�b��
��eN)��O��L{|̫- �C��֗���G�[�6�ad�/�v46��n�/�؅V]������$֟ʦ��u�ȡ�_��o ��+s@g�1�nҗ�}=G�p��<�(o��QbN��\b
�oR���;8��D������s(�j*�Z���j}�����{��qْhz�K�c*���V��lz�p[���v��l�=hG�̈́u�%�/��Y�~s����
}��(���贃T��7��V[`��y��S^�#n�	|N���EH�+��M�& BJ:W�%1�m�}��I�m�$�dݣ�2[�w��O,D{}�}�P,d��Cl7U�F��މ�����d"��+Z5u4 �|ʈ0�dv<�х��p����X���}�S\
�ś��4y�Bʯ1��<�*�f��������O���5���q��G���P�����!v��5�F��PM�V%�����?ӣ�}�|���c��9�D�jXI��G�A`��{�t�ǂ��7i`�%���gM[���` �D��De&���`��^��O;X�s`ۡ] �`<���֥�����j��D9����o�����t8�sWG����'�����%���$����.>-Va�u�i�`\E|���m����-a�fbB������O7�|A�O�&=z��fu��o)����ڌ�VD�q8�&z`~�R��bDf�_�'�Z��2�a��<۳'��lQyt�뽊]3#�эٰI%�l$��&m�.�D+ܝ�����8�q��_.aw���9�j>���c1�x�� �g����҈"�I�3h�E�a	~*�|���0�;���rj�EY��N�
�C_`�G��睌�'��������v�c�)���%�.J@����v�OL�I�Kӈ�XPδu�#nF���?nJ?�a�c5቎�F���5�*�K�{�{����ɒ�Z6YjV�f���}mۖsF��iT�Wv�P�Y[&ͼ�{��?����{�u��
�A�6рcUg͢jǳ�8A�A��&��K��lȊ�"LO|i/oU��lt�����c�r��4�R�k�P���E&�M�����)��l>/���p�w%�ǰ+��aQ��k��k�t��I~6"�n�{�]�}bT�������o��u#����\�cz�
�#_gz���#5Jmݲ���g)!�i�n�Ōb�O'(�8\�W/�?�)v���L�0y�<�Λ$م����ʇ����d宋�q�FP��cbgH)���̪9y�+Fq(:��	���������DH^]T���7C�9��G��L�]�	>u;(�M~f�H�B�{V�[n��qD���K,�Ą˩�U>�#��W��E�Qy����߭��Ct#B��H�s�kJ�-ۙˇ�vR;��ȷ%UP`����J:��U�w�FȻ=�>/nmRTw��#�5ה�gc悹�V�(b�U�p��T> `3�m�z������a�� 
���%5�OZ;w����G�c�d�Sy
ש�]sw=>��=%A�Nv�	b@� ����M����u�+���X*�[m��j�lC�M������|u�H���&�FA�8ߤ���x���S��.�$>d��DCG���vwq�Y{��u�1mQ�5T��C�"fo�,mp�5�Jb��GۍJ��Iw]��lN��?\Etp�p|C-�_H�����ߨn��B.�+��+��x6���:MS;�SР�]�j�'�@r���������P=頄�Q���]M��D�]"ئ�Wd�$"����nX����a�ʅtY݆�L`B�f2�{)̡���*�#��g�y0ݧ.A�F���Ȇ`����^��~'Qp�W�+�9������ީV�0�W�H5�N�����E�N���ٙ�W�7��	&�=43�s��3�u���O�ť]�?vF��
;�Z�{]M���� X�ű��1�������D���l��=�i�a�nG_�M>�R�U����:�D%VH�T�M�S��ra�.� ��iD2�H}İ7T>�pY�ɸX���Z�l]�k_n�0I�'9�+����61e�a�e����`$�Ba�V@����q�g\�dz�k�����=���XO�>E=�_&�<��>���+pC�_��0�Q$
!�|�y�x�#d�ET��'�8n(^d1Q�l�w�!`�C��1& ��MIB������F$jK��l���X�M��|XH���ա�������k�RJ�ƶ*��f�|Un�����Ӟ�C� r�&�]���{����X?��1/�9��oa3���?f��Xvt�}
���'[��wI�FK]N{WRѻ}D�v4���M��S�m�=R-a�Q�����ׯ�i��=G��]�Ⰸ��$f"�RO���&����l��s�9�9����t����_��~�	O@��_�!*">��}�P�z�+�6�Y�6h2P�j����窑}�����PF��H���&��W���r���Pг�&��7N�s��Na��,K���m�&KZ�?d�M>cj�r��.VÖ٦;��=nJ���9�ayz�S=��[L�Nj��1�����?�ݞ�2T�J��G!���X�?��t�e����6��J���!>�s�5���M
�wk���rE�0�k��HiN��f�%���(��+�����9�pպ��`w�Fw$�or�l�H3���-�7F�hv��B�KS�E��*�7 0��Iv+�s�b���3g��������}7¼<���$\`��u��]��ȏ���S�Q������WA��1 �t��i�]3�ŕ���B��V���W�d���b3��6h�w��uv�H@�T�eڹ�V��:�]�g�$�=Y�W�քu��~��o�-vF����Vǐ��f�X�mf�ci<L��y��%X��Gx��#�P<��S5�ߣ�}�퀺��qѿ����V��t�|s�_.�9����Q�=Ö́Z�Oo�-F2DS_����T���1�XN��h�A��l��=$�ć��D]-�+76�œ!�c��������	���on��d�as}�>�p�*�^�_e+�!Q|#�b�6g���ʎC�#�o�� "��Ŧ2�çl���q��w�k	�����ukV���!k2tg���)�h!S}PG��,�[�)��y�[�d� 8��&��^���"�O�c���	J��SNp}���)��;G���1`B�l��Քb������p6� ��(��d�K���ZYQ�x[i\\�?�{��/c��Q>��IR�V���̜>�'FaԶt�pZC��#-+�j�4�{t��.�(f	uB�#�4@DD����@�\�ɭ�BAq}s�E�c���aN�$-�֥˥�
���;��ެ3v�~�+�SkD�҈�$R�C�{��G�_��,G�j����>���B����z���Lt!�󜍒~��ѡ��"���9=�Q������) �����gk(B zA�� ���q��JLڔ��� ;��a�&U�B:���2jC�k.�yb�t�L;�i7Eh�"55��0Ȓ���yf8]���v�
d��^�9W����R���i��C(ܫ�J#���s�u�����jD2~e�y�Q���O2�s� )�����������C�Ğmh�r��<�RU����Eh���a#n��DA_���xȊ����E1K�^�����+ ,f���j#cb^� k)R�ǜ�G.�=ӗȈ�5�UJ:T�k��?H��:�{qA(�8_Ǩ�v`�\� Ot�� ���,K"������ө�{��ב�����Xm�x�:V����و��@*¤�9�$��g�j��z�!�V�4 :�@V,�<G����1�-���߀��k	�CT+�����-�����7#(���]_e(BF����p�c#�|�?E�ę��h\ktr]�a!1]m*A5	oZ���Α0��.4�9�vbds{��v� �U�|��������3$��*�&5���k�~7�;��P��y^�S��V������=݋M7T�V��"c�F�lk�:��M�<��1Oe��^�!����t�ZI���;a�6n��)�#�&6"��~U��{$�L���CP�_�?�F�9��-Z���Ptjd����Q34*��0�qws\WǄ̤W�	� ���B/AX��Ɍ�W���҉�h�L4�����FgU�.��n+�Jc�1w������m���/��"���~��/�Q뙦��V��}B��m� �0��:q7�M��Q��Eh�@a��c���~o��C��R=���F�g��BUǫ��z�lO����Z���������^=H�H����[j��_�fR�%&E���0Z�U<}y��.ABɋ�
^=�`��6k�Ǣ4XՌ�0�Z����/��o�s����Ɵ�����z�>�/7�.�#)�~7�����;?c��k�(W�:����m!����$�-x��d�qȶʝ��OLO�po����#J���NZ��i&{M%Q[[g�����E�9O5�e��$���4����~n���sƧ�;ھ�w�6V���_ӽ�����]�ې}�~�5�\;�Oga O�E���\x3�~�p�6$o���
�{�^?@�+Ie�˃aY�7���Y��  ���t��֝\7��"�z+cvͩ#�&o�7#u����]��,1o�u{�$1[nez̜�������aQV �Vy^�}�8�.I�i���J��>���t��5���^|}�]�I�`�F ��wt�!��W�T�V���`{P�ɭ����©ðy��G�w��6�x>4b,dV�B>)����Z���7��>q��$���ά�\�.@Ĵ����g>Oz�߭Q_Vj.SL�G� ���\u#���ZE�-�Z�Ц	�(��qK�v~)��Z]��(z����].�ad����'���K��Z��C5��m��}��+D��	?�E���8o����$N��~*�	��.j��ˆΏ�� E�`��o2��Ŭ��3�l�����KI\o�J�ux@�"���b7J���)s���ft�T�n�k]�x}��c66*4��ۭ��Έ���U���(��4Ta�\
x2�[B�o�'��d���h.;*�y��p��^�=����������؞�f,��D?���V�ޤ$�;y�i�2���nu �D�B��s()��o�*�I��12�l5C-�Ј�S��j�����/��֟����Ve.�M���q�;���)���U������ea{�{�QO^�
.%H$�]y����+OF��tEG~%�m*����JL�m ���]S�͏Z�E|A-����4���9-˙r8��0���pA=��O�����z�?警+{��fZ
z>�<li�V�fq�p�vO���o��2�	���t>,����c6�^;�?;��O�Ǯ
��j�����<u�ђ�&��LccM0����#���>Y*nw��'`�Y��54���M���q��o��1�W�����F��' A��6}�l�1�������å�Aڹ��U�ΙtH��ݧ��Q"v�!N�%VK)�.��p�N�U0��3��//N��b,_�川NM a��mI���G]�@�bp#7,9Ўp2˪�	�}�	x6�E���D����)yxc�b
u�NQM:���S�F\��
2ԣtYKY�Pe�jw�yR��r����I��٧�[�ͨ�� ��z�_��bE;>�1�-�\�$G9�loX̅i�su/� '�sDE4k�Ȫ	�T���O�s���d�0�P:�����-�ǘ�ss��t����E�"-cb�Tح�"�Z���t�A�m�\��;>�T�2&�! ĻS�B�ekl� zs�F�]��)ބ���h����O�IN4�#>��z�G�(W���O�k�#v�.!'O�)nƯIS��oń����M��=�j�l3��ӟ_<cr�5����7�~9�c�!���n):�~��}O>�ov 
3�Z\��T0u3�������Q�ON�gà-B�U�w";�p�;�{��T;��)8dU���mP9�xJ��7]��&��
� �Nt2�x�X���HȂ����f�;�@E4څ\��j)�MV:�}q7��^�����k�����bh���X�7[?�y8*�  �,ҥ��
��)IX���zeQx��,�AH��K!5����B��	Ϛq���ej�Q����6���O���ٽ�'�H�02Ą��q��kC�/��	/�<�|�[#���P菑m� �!s��l�q�껔�L�2�?�.�z��й?�tE������M(1s�DП�Pū�L�R1�ns��K�EjF�0��o�lEo��A,�̘�W��x�*��������(�bA˳��Z���W��ֿ���zEw�s�h�*ry�,�7��8#�d;��%�yð*�&��I�5�A�ţ��s���������ʱ�L���fg���e���
�]9� �A��u�,b�����\�� aZ���SG�;{Y��Up�I}�{�l6KE{Ĺ�J�^�m�<��������J�c.v�0)��r�<t�z"�\�T��~d*���[�!(ۭ����P�1�H�L��~)?,4��U��It\���ܞZd��j��L�����x�\K=��O��G��d�2=�6u�������mRR�V!r�?����0��z`bp��1��L�f?�K��Klovq�(�V�3�>p0�9`����e��l�1��kO��n�����l����ܕ�u9-��:���O�>x�����2x�м�F�$b�b��M��r٦{?Ǘ��m�Y�T��C� f�ؤֶ�S�R�w�9!�j��������kXk_@:z�?13ܽ�h����eKx1�g�<�ѿ>FN���`��c?�&;��ö�,�ı���8i0U'?���,�'���=X�x�ܶ�T��4uY���)]��K#a�Xo����w�z� �Dzi��rP���
l]�i�˨I�݄5�%r�S�a�:�#�/7MճF�H{�%���y/��U�ݷ|Kf�p�2�?�Ł�U���ك�E:G�� -%_N7B���n�r��E�08���%c������o�@��>u��Xa��lG�x?ޅ��f�e;$Xʕo����{�<.�{�~���ᷥ}o~s���J�,�oE�_�0�/j��m���/�HC"0t�YW�$����N�oJۣR�ϩ�v��1�I�>�B5j\f
+:O������[��Cdr�^�������܍�h,%��Ȗ�N�'�C��r��cX�qk����Y��b2�e�=�@l�QK�1'Z.:���KD�<�:��jܗ������T�-ְ��'�]�-Ӻ�
�a���?$W��$Fq$F�kK��h'-e�o�s9-��=�m�{]�H��_K���O|Ŧ�)2��wFQ������cSp����������7�BLPxH�aq����!���'WB��	H�@�t%�|�o+ϊXE��}L���ud���k˹(H;�MY�.C�7��º3/(XM�ci.�R�'�p�����	H|,�U��F�4㭏��9�'����YB����9��E��� ��
.^��Qyp�D��&��)�U/DÐD�z^�Z��/�[1A 
�-A�J��dcn��aj(G�����bE��A����f��MB]���N
gK�!��;��@ӧ٨v����d@m��D�I�^hW=�ZMA?���D��v�����$�%^�D�/�rr�w$м����_k��y�C����9�cP[�F��d2��ł@�G��mk����/�԰ޖ��>'��2���:��rX�A��u&=3�6���i|�ZN08�?�-�����Yچ���w�n_2�S�J$�vu����7�@j����/�Ti��,}?�v���9)����AS��&�D�T8f���%�^�ٟ�2^GƎV�|%�����~����C����+��|OT�T���FS���!��d���6
	������V �߱�� ��hyi&3��g��Ba3Է��&6�t���3���%���G̅R�]���p(�.�&��p}�{
;��gͲ����[�}уV&���^<��z�̰�s���P�'pV�g}�"׈�'���I� ݿ��xK���:�xm��?���ڒ��I>��HS���H�BE�K���z������%
�t�m��:�vh���|w��)�v����bE�&l�ۤ�|4+ʓ D�l� ����ؠ��+��*mR�GA��z�kڇ�d�n׮���U#!w@&aR8��))��mDu���?��jP~����}H�+�	��5�,�㷂����@X�nCtCV�%�-5�s�Կ��eEqaF��S��̎��FY�
��9U9M9$Wי@W^Ưc
�������(ks��K��Xۍ�:Y%�f��דC�1�%�c�d��)�V��}<h�[�e�Z��Pk|�:Dd�t����]��&�!�L���Lx��e���)��=ݚ	���}��Q:���k��I��u��GY�c|���⹒9�x0!>�z>�=�2U�n�:�CU`�r�K�մ8_��T�xz�	Sc�gR��9�lfR��'G ��9��9O�KRO��2�e��N�����n[�������bE��N�9���2$<����X�ك�uМ�|t3�P+���V��a�����1��_�}$i��y�����䩑��;�Œ��TSwP9���3�����<�X ���mPݤDX��Df�
nh���P����ODS���E5q���lE�v/�W�6`4�k^1���a�e�X&�sPP�28f��?����4Qo�bv�2$&��m{���|�u���i%I'�ވ졦eD�K+�7TݾF~fq�)�)Zc���hN+�<D_b����ڑ��c�d�@�>@P�}���'�y��3�i��o{{���:r�%=,�~�Ez�.�C��7|[̊�(��z�-KE�X���h/�C�b�eM�!���0f������Q|T�S�w�xΞ��	I���2H`�Y���C�_�G-aI��e�x���6��;5
~f�/�X�o�'��k8^R`�7�}�G�ov;v���z<�*iJ���_�$1�Q�¼�Fxŋ�)L��eWג�)Gp���E�p�4�hXR�?��Z���n�����������"��h%�^�Yi;o�ڻ��<�Ӣkx�)N��<��ƣ���>�1��tm���x�P}���@~Ee�qDHEԲ��<3*	9��e�V!�n���� ��,�M�Nf?�;��Lŉ>�C%Ph@fU�=��_��[fW��l\�G��ٶE�����5ND��}wQͿuzqJflF�o�lxK��7�g/C����'wV�Qסs��'&���#��KC~���8ƞ�d�����,i-�._-���� �D�K:��4��އ��U ��o�zK�{��9��G��C;z2$�u��o��gOR���\x�f���}� |lS:$=��*J���q�a �ն���y���^%���EܺCd"')���[�y<��F�ӂ������7w�x;X��X��K�ti-]	��=����p�I�2Im~�y𩌉g�L�jl��Ec?�T}�eǐ��${P�s�����q�B�;�v���v:�791�%uw��"� }�s�W͂�X��#�v4��9t�]3��@���/��0 ϴ�����>T�|��o�Y=ېM�y�xm �%��k�W)SV��x8Q|#|'�ڕ	ι���}>Y�C�o,U��	��`� �n�e�F��ʂ��ؔ��]d�K�Y�f!3�%��C��*��v*j��m��1��wgv�<���ͬ�T���*�y����nu{�ʴ�U�JتUN��j�s~�������0t�Y����o	�G�Q�A�
c%�������!��I��ob��yi�ǚ<�Hm��4�x~{��CSy\Wp�rU�H�@rC�mW�og%�^��J���x��I9�E500���>Ȣk��P;�m���/�D+�:q����l�����D �n
n�J��>�c�ᇥc,��o��U��2R	>h���F(�6A����C�&��Ft\���y�=�否���+���@~�5Ɗ6��6?仲��L��]e)�~�O�/�`��)�ܠ#�J�·sB��M�p�t���8 ��C�2�6�r-E�b<r꽛Cxȏ��K���+����&Y��ߵ]�����3�Me�ͬc� �2��i���]4��Y��V9��K�_�|��r�ˑ�|��=Wi���61��7�dC�Em�s&�L Ա3k*�8���пZ(��eg�[�r�)�1Ǘ�&4cj�D7�	+��\�!�heC��Șz���բ�U�r
}]n�����V�aK�:��Dh�Ҳ&'X��>�J�I-�nЋ{��Ѵɴ��$�u�,�鏴��sn_���8qo����.��+��_�P��2���F��:�u��;�F��q#��H,�h�ا���]J��@������d�g4�����v�R�5i��9n�3"t7J<��8���5�j
�Ѱ.��n/�&QKb0�6�Γ�q;"͑!���xĕ[ⴸ�.@��ݲ�Zol��o�£�t��NX銪@a�����olP�<��.T���M��,���R��	�QV�{�N��E��,��Ȓ�&�@]��C�����_t'H�3#ok�Ū��%ھ�n��|�R��l�Ff8BRsAWM7��$�\��;�]U$a2�`�<�@9$�=��A%U+��%x��e�R�G��qn�	�o5���=��\�tb���c13ں��"Y�pao��ʯ���M>��E�����e)T�#�A��gvW�1aZ@#ndX�m��߬,�/R��w���Ez���-�h���9,�<VP�\b�l���z�����k�՟w��T}�b5$��|�ԧ�(+�0c���^��	����?�*#OL�x�9rW�*�S�K�}��x�3��>�6�1���;��cT�w�w��}W$��*�
���A�p��_)E��s� BG;T�����,�m���sI�j$���➃�T��(m6;��KK����@KA6e cԻ�7��3��-y��	L�1G��y�G��:�/�=���q#�hݻ%�2�l��`M09��5?�LY��^G�]Lh[7���pi(������~����A�r\�[0Y*�����@��C�F�Ů�6Ds-I��6cLNq�b��*��?]<Օդ�
��C`����tA��%��^c�f��T�)��	CIܩ��!Hb�}��v�v��Bg��c�hYn��(5N>.�.�"��{�KC�[k�/��BÓ.������zA�d'!�)�y�l���Κ��޶�Q���]�(�C�׽]k�TR[�EMmh�Đ����<��Íw��g�J���SN��8@�����-QJc_3AV1
�A��Z|��'Z4�~����ɕ�J�X�a� `x���J�,)��7�y����ь�G[���roffŒ8k�?�x��'kfxX�s����ͪƯ�E�K�l��v.-6����U�0l�#!��^_��#�hg|�v�!&$���;u�i^E?�c��u�WD$a��
�Z:x���8#H���XWo�7W�,F��6ˎ�/�ܣ��Ǜ��q?��{� :O�{��^���? ����]���@v�i��^&�<DqO~����G�1��*�x�������Z��-xrC��1#�4/^�_@)v2��-���}����~�w��[z��{22��5sN�L�=*9�8[6�����ѡA�J��!����s{5�]�Κ�C����5b��A��M��Ӷ���c�J�ۘd��[c�=�Li��K��Ƙ��d�y��0TS�3�=p	.�8z�S����nÂ�2��b�J~�/K��F_Ig/2GO-vK���M ����T�>@8�b�%`������pFNA�d&xn�[�0 ��Y��</<���>�r�˔��Q�N5"d_���k�H?R�n�+;�+��ne�2K$�2�ƒS�����;L6�Z~�q��o����3���,H��pbKc-��I��~ �z��U����i�_$C��X�0�N�9�E�vRL�hW�]�̈ y~��k��/V`[zb���R*+D_����"��-�A��c��K��,Y�����
9�n��<�F�����n&�|�A&���s)�Fx&��W-��nQ]��3"b�RnW�d�/�Z�����N�;N�
}L�J���-$!��u]:K��{`�/k�����HI�!�����];��~���'�UQ��E��0k��zH@�^p= Z����$�8c~V���1�-�{��oe��g�Ξ�Pf����K��~�G�۷��]E��y̏��Y��:&+:ne<�#��J�|ԩ{L�"�(�mO- ��L۟9��;�œ��]aN�E�韑�q�cU�v��f��0��&Z��u�������$L���S�F�{��5v��j��U���m���܊C����֪�����LM�/����T\�/��EB^�{s$M!̦��3hloϒ�sBe�\���i'!�m�R�5'���$�͘�\�[����1cD-����{�C�uaN�+�'o���̥W�P>^K�t%�sg�`�(6�Ỷ%r���O�')K�2����@�##���KZ4m�ȵ���8���T%cR�W�L^�/��8���fϱ���qP��9�:W����*)���F����u���-3��u����	�+sNŢx�+'p@�����S-J2$��uKN�������9mG&�\ԣ�C���5�2�9*��}'�X�]�k��&4\n�9t,VB��nc�EB=�~�Ό;���=}`�Թ�߂їR�V����:�	:R��ӆ�V���J�ȯ�f��J�Ľ=Y���M�(�m�Ԟ�l����2���q�V�� ��U�Zw��a^���0dC�=]o�xV�2.@��Ƌ�cmT/�<�0ZA@~9�~�{���X�"��ǚ��$�j!�˒��|�"]�J�8�'��b,�^y��"p��~h�'�>���/�Wԥo�i�i�������e__,M#`a����VR��m�K��0d��i��>q~�F�#�܅�0򳋆z�1�G��.�W��X�SW�����.���=�]�e���<�YF�|�1�%�Aր��ʽٗ���N�� ѭ�%����0'W�­�=6>
�r�`4���j�^f����QZ��-d���h��S	�4ו0�m��Z�r����Yv;������+9�����|�Q0��ɂ���6��(`��(J���Ry:��0�S�>�[��\�:BuC�I�W��� h|2
Y��&G2�> �:�}%����\�)��N�n��44��vX���c�;y&��y^+d]�&���dE���X��d-��BΎم�;��\�7Jɑ�=� ������|������{l�v�ZG�.	����-ױ�%�R�ʵ�K�4��x0h�
�[��'ʓ�?Ӄ�iՁ�e.ݪ���2<=�Z�����',РL0�ML	@Ly�>����犆`8qg�.�r�l���i�y��d�CױA��ˤ�m�Y��3
8�W�t�w�1�5H��L{���
�K���;��~���G]�|��d���MV8P����_����&'
}����EQ.#z�å�6�j���/��m�ixwC��.F��V٪ҭm��Tg���h��*��'��']g��ź����^X��%���3�<��1c�i��xl����eD��*ʌ6R_HO�g*%�ɳ��J�@��H�[����/ J�7(vI|�c���n�MΫ��׻-�o/��]FĮ�h'�I8��M�<���p�(�jSl�Ʀ���ԷC���s��<��R�FO���4��.���w�+��jY��tHǷ��w�PN���qO�)9�;�T���H��;�]+�5�6F�P��ם��`����4ԋ���=2:b���1�ߙ^:�A���D�?��q���:ٵ� �.�W���+=�vAH<��w�❋mڸ�5����ݎ�q$�+�dv�����躄3�e���O��_#�W2�
qE��Ro~܃��o��=�ܭx[^��锿���T9����A� N�kD6�8�Ȏ��`X!�W��̭�!D��p�ь#���E�n�l���:;������v�����P�J�[vx��M_��c�+|��+�|�q�(�R�
�}���/'�9�K�������fVmx���J!��7��`1>�P~�͗\,���Xf��iE@��ʃN*P�*}u曒��+�F��^�w*|ꊐ��*�q[�I[bX��[����h�qQ��V�K�>���of����L(��$j��"g7�_"�R�������pڬa����~/�x��� WK��}�q�HG�Su���[6j�Ӫ΄k��d�R*���H|������J��]7oi�7��h�7kH�����9}O��@'�%6�̞Ǡ5�K{��;Y�14�rX���������C��7"Y*�7�:W��3��O {���k+���/o/P^�r���q���������p1�u��p.4ߌklj��������}Nc�V����?{�9:d��X������=U���a,d�^�jd}����\`�� ����8�{z
�Tyc픛��!M��%��h (dс)y���9yӌ��������~���|ي)H��RXq�k�A识�oq�����ϻ?�>j�?�ɛ�V/2�(x$�(I��,/�AΒ���������v��7���֪�"s�={I�hX�Jyg���a{p�Vm����P�ڔz��hTWV.�cb�{�к�s�(���ù�9���>IֻaU�l�P�<��.-���/oj<��u����Z�zW5���mE!��x�DOD6IQ�� ��� ��k%��2�i�:�M��6���q';�X#���?j_p��8�zJ��ݲq�"l�*�Oܟ�,���J���/�G���OW��欌N����o�\֝�M�%I�`�E�y'J���NI��ﷅ�]}�����OO�6�1��վ�T��E�q�|�0V� >}E���k�y��L7���9�6ڧ���u��������H���D�C��>k�6�ZY�G�x*A�`��`�{_-j��5s��N��HKQs��cK��P��6~Q/^��2&�͋��_ԗ�3���&H�Ps�3E��x-�#X�&!�d���[��-nri;:B�Y]%nM�4� {�(�hj�q����P��T�S/b慒v����Y8X�w�On5V�{x�1��K�X����Hc��P�՘������D��j=��{l'����q�����i�|���u��`l;�;�H�
�^*,�ݿI��V
�'�u�M.��\3L��҈;G���)��k	�⊿�Q�D9��3��5���� �����l珣�E�(�FQs���|���^Cp���vi'�& "b�.6NF��+b`�K��������.	���5��H�y�6�K�*��4��,����gM�\m-�)-Č��	����C��Թ_�����P� E�C�Kz�&=�@o�����d�- Lo���^��(?����>���>+u=�Q�ё���ޟ�h$����<�G��G��{�ߛ���R�1+u�y����!��o�&՛\���� h�mZx�� ��I�mФR��U�Mb�U&�3'�#F��v�����A:�����$�������0�3L���!$ҩ��Ua���<
�B�&����2y����7?z�5<G����p1��AI��y��ّj�(���9;B^��z���)���N���8&*Dj���/oE+�>�� 3l��[��ɔ���7jl{ԭ�':�I{�V죭C�-����5��+6}i�qǚr�\E�s����7V!�4��B�m��g�ּ%&He�AU��Q����<&��_��E9ks�^�,�����>��С�8��:��Z+1T�p�!�Y�t`4[y�?��k�I�H<gr�$�֬4�վ��gl�	��9a��/2�����WLX�����`2T�D�g�{ݶш��&��˃r��Ȗ{����k�LS�#а��n�k1�
�R�� �k�%�d�Ո3���F@6p�~n�[G^�
�P�Bqp-c�@��u�
3�AݱGZ=�#�=�W��G�cHÚ�:#�"H�K�&d�a���ڬ��x@��4����ć���4$��� �}�Zt�\+��;A�\��j�~�;�/��0c��-�%����׹������}�UV�Z#��2�ja�D��Jx�廸�0�]���ȱ�۰�?ZBȫ�gp/6s��f��w
��&g^9B�]�#7W��O�,¨����6��I2 	���$~W��te?Z�5ڛ�R(��4�%���G�N�n���c�����1���.:jT[}��\�;ܐ�x��d��#�?�'a���d�J�y�Z �-�B������{�g���bB�!��@G�7�XC�ƍ�]��<�x�Hh��ц�p�Э0����N�6S�#� !~��T@�"�%c�=Ӵ�R���虧{�\���ѠZ177�}X�������-�Z{���3,��S_�Ku~��Oz�����,��I��R���7%$sU���8gKq"�3M�*$���bʯ��'�$��ݙ6�Y�������~�q�QtE�.�����u�B02ztj�v�ⷷ�3�w���1{
,}�� ����V�8��m6�Tu�ն�q_�L���'��b�I����;(�T������h��M �����Ki��j12�Zj�sC�����M�G&y�C��Mw,]��V�d�o_~DG&f��|�l7fM����������x_)�|A�rF�kz=\}PVE�."drڦD�����Q�MA����A�N�|L;�혜�� ��8�Xh�xW=�Rƚy� �l?�o�)�u88���Fe�>��l�l����Z�ۨz��*�d�e	5��=1��� 8��>�`�[�۫���	/fݏ�䖠��r��sl~k��5��Uִ�79RW�ܠ�w�Q{?�L�*��D�� �]�
k�Q`���m���c���:�ev��Mz���(���*I�0������;�ȐbN���]����b��t
�(7��Bg[�����k1yL �[~��#L�M2c���d���� �m���A�q=bi���+��?�5����m׍^}�ݖ�0o�vher@Lw�q��A
'I'�{w�_�b$&o��۞#+�ߪӧ�a��]���n��m��� ﳯ(��/�^4��9(�Y@U��Oƺ�x��`LB�J�=�ٱZj%��$A	R���</����1��ݵ���������̀�o��~fv�Іs�˿�q��G�ׁ�d�B&�N�3�x��q�������$W9rpo��	�����U9�="\���5�� G������v�oX��>�gBA���#238Dx`��>G��ŀ���^��+-��ȃVy���b�`��	�N�I2[���$�a_������p��g�Ԛ�G֧b�;C��~�S-%k�锤+�>�p�r���N���>.d9�E�j�3&?��.��F(�#@���S�ya�{�T��_E�^ĂZ�?9���j���K+���\��,�@�눩���.�[�^��I�=�7,�)ɩ���:�\�6Lo�<\{m�!���ز͢��2'�T{9�հ��)�"\aYV_t���Iq���D���jv�S'���$� 06>���J1-H&����[�J��6?�F۝�E�SN�Q!�|c�h-81pS�Z��G>�{�0I��~�B��h&�"�p|��Yd�ۑ����8��Զ.+�l:��z\޾��9�����
�ݽ����E���dECQ�Fgx�',�?c�"?���m���:��w���*��^B��V���&�������}9�4���(�iL��k���Ӯ�n�Eh�.-3��t�X�[Df�"�G%�U�k�LA�A�ǿ���U���V�0Y�a��)Mm �ܩ�(v�PM��c.٤4���U1Us���Ęx�2]i1�9¯+87�b%g�.�z�=3�ӆ8b⦩N�Jܳ��S_�IZD��#j��?bV#�f��{�0�~^��׾ʳ��bţ����8C3�W��mo��rC�P�YF̫�j��M���2!	o���$���w~C���b���u���䊝�s�<8Ȣ��P��h�d-p��o˾E�!�k���+�_wd�T}Zw=n�c"p������=�`Ԃx}	�+Z�O�G��4+(m��87����Y��_a�����4�Z�D6���?a�D���۪����BȳBp/��P�ԙ�<���^-�z�����Bi+��1G���~��Һ��I�����������H��EU�����5��7�� �鮫oL�Me7��;�~���8�zV
l���ت����2��1Ov�{���\J�)m���X�+f��CV{E�EM*�65$�cʂcԗd�щ���nA�(KV��)$�Scdʔ�y��9����H��C�ِz��B�`���@-�|g&="9*��y�+��)8bƗs���1.5Vl�1�2%�դ�9��K~#��!��R��k�+�B����=Zc�U4�;DP�:�SE���ۢb`3��\wq6�>=k1�FM�� �8K���r�`�t3�Ixn�J�ds3V�E0�tL�*�+l��0�3~�kݼYm;������2����6�@�����|r)>{)��0}�:.$�/I:ř��q�d�4�^�cư@���3k�im���)�[�Uп�Y���F4�;]�j�`_�+��j���li��%Y;�����$�'����He��0��+\܈A��2h	i��xv����a;ϓ=ٙQ��s��:ƓE�ʈ�,���Uv��xdr��w���fK�������$ɢ}=�oR�xX�|d��O���1�y;E�`�Cjΐg�P%���,��׫�s�]�?d.Lf�m)O��\�+u�G���^v�zG�㌭��O��z�`<u�=��)�ۯ�����p$MNI��� ��i�{��9Ԗ䘇خ�9�ka��8�cJ/�,|����|�p�X�$G���4 *��[���qƊ��;��Z�k�aU��xxt���8���>�[����/i~�z�q��~�up���r9W��� �D@/��`�"��l,���R���r�뇟� %P��s[��w0�)����y�jh����,fq�[��M�Z�>`X�y}=�.e�[�U�4���N����H�¼Gc�W<"��dH\H]3s�}LPuϭ�t4�Mg'�� ��}`������{�]�3��B9H�%<�)���\z���w��#{��w�XVt%�S���L�6r�/
v_~ͺ*���yi�����\+a��ɶ�\�(��t��ڮLH�k2;B篴����d��~�T���6��lTYeb�2?�\�CG5i�s�C4��NwOw����Υ���$�����m��`����a�lJf_�kh�Ab�����=�eP�� �eċ�s./`�O}}b��͢�Y��@�?�����!���|k����T(��شF�R�_��%v���̻��W��m�^�W��;�)W��c<!��z�b/���L�
���~Acr��1���o��+��5��l�@�,��]�Yw�@/dۢ�֧������}Zk8����5��_�`�-��4�铮����?�}���h@C���3M6���VAxο�B�����`ݬWh�EP�d!PU.�Fĵ���?�1J U,�ƙk����>��"A��5�C��K��B�����l#�Z+��E�H�����޳�[+-ꍷ{L�=ó؍khFm�ΞKH���9*��˟s$L�v�֩Ng���j�� ��~H!<]R�ԕk�zc$�����;�ܪ�}/�$�J�G���m���
r��P�qF%{K�H[i�=9)Hz-ǟ��g�CIh��b6K��w'O�Gm�1%,��	��'�P�^Mp"�z���b⢆"?�hŚ�k�&��%f�:���DPyR�
̧��h�g�Q���=�X,�
����L��"��ߙ�K�)�?s.��zw���-�~���E5Аqځ��qx�X�P�����Hb�7�JZ�qL盛�h��aP���)L����x��m�12l���=T2�[=��� Q����`0w�UmVÿW��n��E3�q���}�aݯ&A�޸n�n����k5����{6�����nad����d/O^��c��D&��%�}�7?���`W/�s]���:�	Rrt��� '�(1v�@�[nGe���)�,�(i���aG�wo!��u!�V#�Yە���Hy�$���~���-��s��˦dW˫nk�;_:��)��G��d��ɶ�E��<����ERm7a�����P�٪�#�J]�ǸE�|��?��tkh]�i&�'0���̈́�����vĪ���,��-����^�B0}�<�c�N̾�c�p]��q�w�&��/����+-��ߛ���ë� '@b�{e�O� �3��s}�י�tR`ܡf G���y��� �Ŷ9/��J�Ǫ6�@]u�w��I�X!ȶ�:�N��dm��T�x�1����P'��}^hZ�o��9����ۀ�NFiR���Z�թ�ʒPig���Ӑ'���YH�]pЙS� ��U[�e��mf�cB�1C0��5�5O�{CG�p��0�y�:�_y�|t��xtP�&���4WX|!��,w!\�� ��R'�6��NA��O<����Dm�P�'���/w���FQIm�Xv�Y�҅�:Lb�oˡ~E�\��V�F����95�,�v�Ȼ�l?���t��}oi
��Ֆ���%�r�E�7XTMF'�r8����7�l i;'8qH�Ո�����y��V����`��Ί�Z��f�!0O4q}Jt���S�0���W�;�ff-�-��@;\g-�)��6�-�����`�}�2M\T���"�<�OYe-�h�ΰ&1E=�b�������ҿ�ϝ�ad���P�Sgc��B�do}����a�i�ӎ�F��a
0��HIܕR�����67�� ���I26"�B� Z�b�M���{�Ǉi���*f�?G�W�.>IH��Bv[�������:�ް:
��m烝�u�R�{�i#Z����#�t<�d��� }uSAh��v{�G�5�7��S�?���]�8��� d�[Q�!����v�:z�Z1~xNW�F�>�jC�!P���?�3��1%�;^3.��`N�I0c�^����݀����UCl�����9���L柑�yO�W}���y2O�=< %R�	��a�2�o�Z��{)����x�0�/mt�L5ؾ9�^���0�^{^�������J�v�Ĕ�f�(�o�N��*��f�؂�]@�P`b����9db䖄��7�9Pв�ϑ��~?��QQ���a�<����by �C�<h����
t�ptzƯ��A�:D��J׫|]�[W���7:�L��Or��!�9������q���X.t9v�QӅ���?}�/��䣸
�)�4A�%e�'& ~�;�t��eԘ�~��_h]G�8h�c�1�A-�
6�@�5�eO�c�HgW6��R�"�:+���G��cw�2��KR��JS7��F(w��K�-� ������ۿ�rR��EE.v��
���/����/C(} ܲ>�(D��w�upJ����.+_�9)[Q�sVB��q���ކw��[L�$g��q�&��i�GT��ך�$U�f@���G�p�_�ݳ�TZI��� �,^κ��k���ޙ������P~7��fVŐ�֌[�U��4��$�\�Id��;��A�Q����b3Y1�p�{|�5jM�T�<\�l��N\Vtxu�~%���k�_A�����'-��ȗx��\�$�څ�?�d|n& w�
&��8�����['����q`a�_���.��5�/@*\�ࠢ�kTo�q$�	����C�$�������z��~� i�mRfR�ŋ�ʲ���Ns��f�<��1����wW���1$�\�����{� z�bSOl�(�VB���9S!"��!�����u�My�:t(��F�CRpP��Y�=<�\*����`f���_���\]��Tv�Ȥ%����W�ou��oc�18�+P�m��1*�{�&*�� O�Jw��E�����w�N����^�m2z��(��x�I��7j��C]��5��([e���8�|u�\�ub�BirN��7et�ďV]�2z@�~�Lpci���s�b@���2i�e��Du����t�f�d���Zy�A��Ow_T~n�7:$��2���#j���I@�"=Ʀ�]`Eu4삕�!���)X���OH�ՍS�T#D���q{��p�RTL�:e4�w��9�Vƃ:_f�d����.m*Y�_�#�8�
�ڧ��Q�^gM�y�kqO��<�x�4;���{�3bsM�}N�T��f�%�amٲ;��2FG�#��B�yTQ��E�ߛ�Z��2�7��/}q��Iݭ-�8��=�R�'��O�T'0��IP�u�t���}BO�	�`Ӑ��(,�@��b��0UBU�fq��ZD�~�Q#�O�b���x��w�i��*]�m��_կ<�z�E�k\�5,[5�Rw�f<N)=�O��8zd����ܞ�̹BW���E�C^V9s��a4ɭ��QM+��-���Z�V��*	�\Y��ɽ�Y�S�:X��L��~�}�&����`�ѮѴ�1�ũ�h�N4	~����$͟�`�J6L 0�!Ä�Fq�<1#��!!6X�le#on���`)�WZ2� E6R�<ۊ��L�ľ�z��_"�Z�;��I+�����)d��g��ڼt���]P9��iƊ�hȰWސ2,�_�⾓���eR0+Ip�T�ā��Vu<S�{��fDv{h����u�Ґ�)�r���A!E��L��r~�L�b����%�VE��+vs�\RNI\�%/_F�x�e���U��I���n�SZ·*!�"ڹBU�;3hiq�Գv{�I�?�:G"OT�G�%�Y�
��ToK}�_ -� �� g��'��"�x����������M�=I@\$���O��^�9MZqkꥪ��?���o���t�J�����ː�A;��n�P����/_�e��i9�"�V{k�Т*�� ��2��)v�R��&�[x"è��Y�iWQ�vN�F���f�q��k}RB�-T(yz1qB�4ZԧV[����Ȁ��i�a�!怋D[�2��`�adp�%8���Zq��!b㰩� �4L],���R,ҭt�K�eXٗ㤕��$Y����"~)=�M�!���1^����z ��"������=����#�tVo�KC�x�:�F��$�s�Q�H��ƽ�q7=�C� dO��'� �_����-�es|�H��Ψ�W�^�[�T�Q
���KpYA�Z#ʱ���Q��J����<${����h��$�NX��E��k����fa8r%�T�j�@�𘐡;N��7�

����[�+>�t�S�Ӭ<� �2��[���gQ�쉆d����Zwݴ�8��{Oւ�oA�_������S1��;�v��m,�@ Y��#�]�y������D-�	�"$I��/��,w�9<;G����c�^wV𲪢=?������ӽ����!�j����׌�r��˥7	h���ek�������@�J[�}8�^","}-��h7j�h[�՜��C}.�.K�\:�8�׾+O|G&�N�Y��y���/�0���W�S�XR�,]��G%׋v��G4�0Y�*��V&�/��y"d;��GU8f���12�Va����㦥�7�{w���>A1@rT��o�Ez�)����@�1X�J�99=�����
kcx?�mh"�y�风�B�ǀ%��.Gs[�:��:�jz���t�9}�u�σ���.Ke���~�jцGiݖ�:
��)s��U�h~�vݜLem���,%}�zUƼ^��"a�?A�9���,׾���c@"=!��{|8�C e���� Vi��]Ϙ�Pi����qߙ9D��sP�O}E�F�{���,%yu�����v�3�OQ/���qi�amf���&��j�e��B�("����`�n*���~H���1m�*a!��.��%]��b�q��٫Ya5�$���np
R��#��CjéjD��ӯ��ᕡ�R��W.qXI$+a�'IHI��/��ފ��75<����!#��S'4�60��J�X���n�䷷*�"���1s1��Mx�]Xܿ�M���I� ��#�Z��j�Ƛ-����X���X;_���2r�^Ab�mF����MX"w҆��k�r^E��9�Y�zT�tKE��������'=��m�zJc�k�d�j������)Z�#~[��k}� Mon�j��1�۠>p�l>b����5����ౄ%��wض��@�
���k�2�q�ڦ��z���v���}��L�ƛ���_�%���r��"SD��ds����s�t$B��Q��Q[)%"d�ń�ʵ��a�I�ߦ��9CGM:@���f��Q���߃>k�(̭<W�p�q��9��k߲��;��CS�F���y�Aic��~���K�g��d7f~��
��2] �R�AV�.3�6�|kg���s��-s���&n8��{�Z�⇠"��s���G.�op� ���d�y�[Ǣ���nȋ(���O��T\��f�s�`B��Z�c�t�j��*��2��[�ۗ���*�s����E���5���wH���i���u�wj#���M!�BL#������I���v��tܝ�*<=�Uٵ��g�]J�9�W@tp9ka�x����ǉ)4Eh(�Ѡ���s
/������E��u7L�"\���0SyE6�8j��vAh���/yնp��:�O���հ׍�		9�ֿP��
:qby=�/�9rKQ��+��xOΈ�>䑛6)W���78�m�5)<���y�[?��&�zl�MS����$�ɲ8��@�?m�a�au��>%4�9��]�)�bɖAJH8�&��/ySd�Mx	o�)����C(��~}�?��9�
��O<Z^_+���*�ʤp�n3
k�Ƽ�Gr��^(zs�p�I���Y������G	�h&&N���6�UIU�a0��|�1���#��;���:�p��x�R�y�I��!���?��q��;R��?�P�iɇ�C��bb� (��U�����03ԭe�0<G��������E��hO�孔�W��GoQl�B.���9~�q��\QcF�3�[30�uZx˿�9��+,=W�cׯ���	qCp:[[���瘠L�VG
/�G�,��C�ֺ��|�C�������}i���7�^�#��m/�r|o�c�vxv�琑�J�~2\���� Î�R��Ra#Gڮ$���$��"Ζ�K:"R_w��d�j��Xn�:@����ʿ��	FE+Xd)����Q���B���.�W�g���df9�������;��h�RF�ھJ�_;��5Rr�T�� �{o���$_���^sϛ����Ic�5K����s�/ݕ[�������(�cK�K%�ڦ��t4��٨�LnB����!:W+%����:����f�d�I` ��h����0f g��_'υ����1��@�Ǳ�$W���4����3ӱ�;�' ��n��qU�+��	�r�hy�6ԉ�k'�)ߺ6��p�	C�B���*�B�����>a�(˚���H<�_�ǩ���g�����L���Z�!v������P���аh$5�(���'����+}i�(<_�&kxˆ�;ؑ��^>������^��K>e� ����w�/�#a���U���l)L�0�ҡ��'�[�vmZ�i�� �݌%1F�J+�T��������X���%O��E�E,]��{}av�W���u�#�ynDĳkD���O���sȚ�f�Y�T��c��	�m����2��)�u��������z�ffu�!k�U�]sk���75s��r�ýF�&SF�1�C�T�dhʼU��X�J�T�kC���>{�+�:����Hj�)�%�)�S���{c3��x�6ߎ��z��\g	�q�V��
Ī��	�{��wc�z?9`���G�&o�;�ϋ<���P]qZֻ�ʬ~�}ƇM���!�5�[K��+�˄f�~�xG�h�G,L ʊ��� ��U��p�5�V���<ґ^�o�����ފ��fI�]���T��^в�^:@%sqV�.��4A&E|D��)��o���S���u���?�&�_�uS�q��:\K`�����I�ޥ{����O�6�Lz;$b����[����Eی�M��6`a3��{��ް�W�����/�񝔲B�t*J���I���1g�Yi�c�HQ��P���I����0e��ӑy�����g�0(����4�H����o9o�t�n0���~~Rn7��߁��ǝgN6�wpWdOS ��y�B��=�!�ï�F���#���� �bP^�!�E	�����8hw˗6���n����ƽ�>�Ss~�]�U/�?�oY��0[�lŁƵ��sd�7���,'Rz��_����h@���s�u3²U�a�?�#p�髧���evC����Ʋ�-T�Ò4��Y���[��Xqgt&��|#*��߼g՟��UTq�쏎��EK|�ݒ�p6��G�F�/(HTsD�Q-����r%��_Pݨ�4���M��Xp<����*�<�^��kN�R#���ݕ³\�@��.���o�M6�Ew"Q�(z��L�˜��� ����v_Q�Wj���C1��U356g��v,��2�g��8�Δ�#��!f~#�_��.�r����FyS�b(�R�̻���>%-x�f�M����0���~�V��/6��*j���T!m�����,>�1D�����b�4��
��h��%��c���;E���t����Ă���� ۚ��F�x�,M�W����ql.����o���F���&�����<ɪ�����<��ܟ2n:�%�0鄎�{`D��yO@�[>IZ�yf��򆆏�F��NT[x�V����C�qE���R#�ڏ8�CveX��9��F����C�<��cKLǽT�o���܉�N���K�'˵���KL���!r�䘑ף@�V�fi�(�G)�xd�L�:d���(ug�΁u'v�i�wbǛ�Ej`&r� ��4����p�HL=��g��X<�ʴ�Ǟ����Ű6���Ěy[����u���E#'2���X&T��@��z/�@��$�#��;�� ��в6\)�o� �?N!Q��|QW~����I͝5Ya#�?[8�P�x�~c�?6u�=E��K�y�	-��گ9R��H��� �¡%�5��u���N�5q��Cf���oU�F
N��5yL�,��6>Q��3q5P*�qoR�r��u�� ݵZ7vv��}1��F_�y�8C�P���.<y��Ŕr�m�_����ΰ�5���)��Zʦ�3�\{�<%�Y�L�������]�Os�R�����7M"�xҞ����)NU}-F�T�E�C/ԃ�8�։��#��f�Q��Q�i�� �Ěd��D5��L�a��>R�F���v��{	�H�l��	��^4U�m��>d�S�6���-ܳ�s��g�yߕ�4�*�<�I��7ەnpe7M����"�q���Ű3��sa�ɬG8&���C�L�w���.X
��o���r�z����gW�9�#���Pg�t@%��(�����&;�e�ƶWC����<W�4��*��q�;p�D�o��Rq �J�����w�Z h@q���'\�?M_Kn�1y=��H7�_���צ�Ѿ���|��~�wή-��!࿄8��� :o��a�t��L�����G��U`����B����� �reT��#v������蒭˝�-�&԰�Tʤ8gB9��U���}TR�@�k�<8`�vEܼ��I�E��PV�M8`��t@
��W*����Gx��zA��EG�Qʁ�t�5R��?�O5I�+Gwp�Y���w؏��5���!0��I��a=K<8�3$�'|:Y�n��a����Vu�+ŷ�,�%��R� b$����Ćf0�i� &�=������X3\{d?{T�9K3���#�|�8m�Ɠ���1x���V����ߜ9��hB��	���8�O ��o�e��
�^��ۼ�P���������+/_m��;ӂe{ox�%�Q~4��w��g�2y*Ck��ۙ���f�vNvxvC�dz;�tY�U�7 LJ�ßd:��k�x�{AR<?��y���|0X�K�*�k9~P����m���ɺ�\�~qF�֟\t�h�}�mŏ�F��F�-4S��G���&!���tÈn��"�V^D>-�Z��b�G�,�Npr�c��X�Q��ߋv�Q��@��s�ڨ����Na�d�,7�#=��7���)iX���3$ƻ=:�������5,g�����Zx���%t�� ��M�8��B��Fd5�h�$}С���Z|��Gk���	և\W�\Rׅ�/�[	@����z����~ca��x:�m�;��mj�:���p�A9���Ft`L3�=K���<3J�
���.	�'�I���+����T��9|���!������(��M��1�g���#2	Zv9�"y�$C���n�H�;/M:}˝3q�K����䖃
�KV��?g��|�2��|����j����7�iSD��).S�e^B���U�*P��m�DW�Q-;׵�#�vݷ��I,\Z�ΰ3`9�A�WϺ�\���2k��%���B�D�Gj�q�7r���G%����<��6R��wy	�$C`�Fj��릢����K1����t�0S�*@����\�s斦�G�Qy�s�̖HN��j9��/<�5�.�[�G�Ӟ-s�����Ћ7�E��z�u�3ĝ}Bnk.������6�wa�!��aI�KnhR����ᄩZ������Z�gJ6��~e�y��ƴ4	��m�����3ha��Fi�\}톳7[�_;��[�ԑ�ȥٚ��`�B"���jL,G�(��m�`:��sMr,�(ʀ�� �A�{�5��v���u���j�@�Q����+&4R$�Y�d�i[p�1k�>P7��f�U�e��>����GY[���������XuXp.Re�b�$^�L�2R��i�9h��Ű3� ��l��F�q|��6$~<s�L���y�5p�9�;p�\�G�Jm$	{\#Œu���Tb��h�� �b%N6�Ǧ��S�����H�X[q�./��J���v ~��n��N�Ƴ��m�L���F�.��&Ċ5$�Ӫ'�J��X�S�dk�Ivh�ty}F�%���rf��E;��A&r��B��*���dPsɾМQ̛4���V;>����z�0<�(���i�`/a��ވz)�!����C�(�Q�Ƃˊ@\�5Ř�þI=�R�"h�l��R�s����6�&,St�/�l���P�{�d��&�9���h���[Ľuɿ	�z;�6��qrEG�u��q��ė9C�E��1%9+P�HUp�#L�'�p�5A�A�"�=�}���v�d�E��m�� X������E^�b}�Ȉ4"B�1�{���@ �<%����չ?�SA��I��������3����F�S�R��'�U�dA�x�h�E�/�v@����J��Ȗ�L:��6�r%�3�` ���*�����wI���\ؒy6q��r%���Sr(OMR�:��'EI�<&�Ӊ;r�����4�Dt�8Q��'�LK%�rE�+�����CE�v�����HOH�-��~��Z)W
��8ֳ���ݐ�-�=<g���p��t��:�*��Ii��#��Η�u��oYrF�OCn��PFU��:��2�̇�*�Av�����@�EH5G&�[��9��L>L�fG�s�@��2�T��2����0�ҵ�A/��ն��o�v��!7�&��n:�x�ް�*�@�N6�&^$���L�
2s�yPf�5(�D��B�u�C?d[��DpQ��#+�*�2TRÀ��%%aY�É�v��Յ#�`E>��C1hX��}'���G&���%;����
]�7��1����H]�kj)T�ʾ!\ؑBj4��}\����B{��j������D�����J�ö��
E	$H���/��w�m�;��*�{i�{�[kQ��r�z�6�8d�� !���M�y��N�'�d�ۆ�#	BZ`�.W��\��+�̭X3Kb��\��=I�=���hL ����@��)�+�2�7��Dd4◤]�~A�#r�g-�H"O�{��<�~�Zz���WZw{�f9Ƙ��=�g�C�ލ�^?����o�jcH�E\O���`�е�d	�����W����<��;�o`r�^�W��}d��n�1�v�0�%q��*��A0G���j���W@6W�XnQ�����.�zf� 7�z����,�,�`��`�U =2��xj_d��8Az;�3�rbM����<� �=9M������?�؏�g��%.3@9ņ���QT���D���3����+����*��,+5j3�I�h�L2�N���P���tS�+��^n����Ku|��al�4��k��u�8�hMZ��6���q%����Am�] �V<ꗅ��O���1����|n�ja| <�A�SZ)e����4n�v������ zI�r'G:�g���(4������Xl�`�5�5v^0�����Ds����T�!,�Ůn�����d� /Y�xv)`�>Q��z�����E����j����_%����"��R<qo����9��"���M�s:?`j�O�H�;o\�q�E7n����C��(У;(�c�)��d��)���QF�����SHܨ�@}+~��O�S�d��wnzw��mB���S���J� �,#��:��c0������溰x:�
���!b>7�U]B�S�Փ�D��G��C�lI"^��ޮc�"����� w�I�'	��-��U(�%@.5ي�m4y5NAVh�X/�]��S�@	�c���c�������������[FL��t��'������O���ZBe`b�lڙZ�Ht�s%�e�����5*]�$$��z˖ʟ{��
��)��щ�0@�E�8x[���Q��D���\.^\�6;6��K���Ѩ���i���*/��~H�z:#�3;(�4�b��A������[�����cߡ�	,^c���*����YR�m�D ^�&xgA�2}`U)ڿ/�`�M�A��P{��FΟ��WS��h�D\g��x��^�5[�~��o,��S��U����F�Ӷ�?H~p����8��}K	VY�]�0�D�G]A�M݀}3�^b�,����[�l��cm:�:~Bu�l�!�=�"qې�y�>~�~�Hjp
��%H����Uv1ʒ�	Hx�G��T_��^%����t|����ߖ�����:���m���j������Vo^�n9Е,�I��b�[�V+$D���Q��Z�����9cQ.�כ�H��>����0�S(uy��Ȏ�p�n�V�T<��d�o�$��knDN<ɔE�	6�/����I;$��F/�z[��<T��Mj���-wY9��*@f�(k� ����x�WG�aK�cu��m	��ra7 ��J�uݓOy����oc���knk�o�ˁ�h�*�B<rΫ��W���y<B}p.��ο��?�՗��t�u!S6g[����?�����b��1�����|�'7�غ	I[�	�(O����0��qxa�vX��xX���m�#<׷� ��?�L3��Fx�g��Y�:�"\c�'&_�s�Q��ɮ�3�K>�yg�F��mڂ]�Ǆ��L��7�+$'aa{ո���8D�l�K|�g��n������4f�Z=˅�,�~�g�,O�it�
$Z�	@��G�n	�]��տC�aj:�KWFM�B�����G��$�
� <Z����s��/��-.ycu�U���I��;��9蠧������+s7o[Y �&�� Y���ú�4����6�1����pXz�ȉ�������PR�t@�,����>^�e���H���P�>t��T�9�"Ô�>��G� �m7Rm���蹐z�}�/�:�Ds7���MCmf��h��w2 &���� ��RU�ς/�-Ё5�\Jt=����`)vl�Ƴ�J+D�>��'8��[�����Kt�j�J���di�7��N���AD���󱰞 y�SOs�ו��L�m��Pcp5ȶ<�6P���@!˪Н�nd��O�ҧ�,cn�K�~��9r;u�^9�N���,󮟄ӄ��%��\)k����x9^��ۏ�6�A��6��6� ���0��� ����:]�D���;$yt��L�H�o,���W�: ޸¨6���a�SG[\����S"������p�z`B۶i�����ݲ]�_��Rb�A�YO��Fz
�xj���5��l��{~��>˦~��Nec���%h��YNW$�5��E	�Bͮ�1�v��3w�޶6�E���c=�
!K�F�R 1�)a��v�B ���4茦k����(�q7Ĵц���'��ƞY\̠�	Zp{��.]%~)�n��S�q���h�CRҜ7���6z�nG�T��e�4�E��I��ѭZ���4��,��e͕-4�H��,����[��b��.rzkĨ��"��.^�������/~!o��-t��=L�­�	WNYW�x+1(�#��C�Vejb����> ���͑��(���
��$)^0I��ٛ��V���t!�G�f���;���ظU��P��F�E�W���G���)�$��zN���0�:�5�#��1��@j���^}U�`&��DV9Z�í��� 4�R��EX�w�!~%N�;���xQ�\}$9$�[E-�8��?o?�H�g�8x���;p���:��@v]6G4��|o��a%ܡ�ln�T�G8f&8҇(=��a�	�J��B' w��Y�Pa���n��G�u"6:��dA�9E��3�����&���n��4�.�I��Ήa� s	��Y`Ro���gC�gI���a�4�;'w,d��l��$���]�aD����n�e#�>�k~؈H���2�R����{$ѓ��$#�qms��o�?Һ[W<����ŷO>ڐ�v�d�x4w��ӷ�D՚�3C�u�Yr�a>��G�d#=�0�)���۞/|-`�0:�y��9�y�ʋ7�� �q��Mt]��q�\��I�4�H(6�ԔOsu��>�9"&KD�2[ �'��3{���ɔ{���=��1P?9�8���ܝ��P��y~^��"A�����4s�a%�y�cӮE�Nj��/q���~4'�Qr��\D�ͧhU��4�Q���
��@|���z����x��=�;����������Dv^�.b�����+k<�R����h��?^F�[Z�{�M��}�>Z�2Nc�������y����⍡,��Z�Z)7��e=�D�*�U�A~n�K��|�rm��m6sZ�yo�b���k����$|M�u��2˽���Dy��B�4���wF���PUHf��v�R5��:�bʳ���=V�K]��.�1��\�*��$H�0�3��W�1,��`[J1�ɥÇa�B ��DR���b��
�ƣ��ŵ���ՒZ�a
��g���!���,P��B�LNi�V4h�r�k�����8'L1��x,�쯚�d�*��q�Eۍ��֤a������^��[Е#8}cD���T��/�čX,f&=�=?�g���)��gknT�qG�Y��pX��]��>�"�]:�:a����?����Et]k��LH�{Olj����pL�e�O�L����=��-Hj(��4:��l.t�%�RL�j@� ڇw�fRX5h��7�I6�=��"%�u�a��VV�[ �*4��$���9��q��7����fl¼N��1F�5�,nUJDեhy�Hn�&}�KE|��?��y&u�uћ��pݣ,~�u4g�MQ�ϲ��Eg޼u�'<���kބ�k����H���/��P&��X�� �<\Q��X%�`���q��ˠ ���"�?4�����+~��tp���(ƥڹ���w!V"��6�h���ǿ,V�c������/��E0��k1J�X��� �B�)˿[�|P�4��Mg���̧z��_���\�3%e��	��᪵~39ޔ�㦼6+F#y!b����76���]3% ��N�^���Zm�d��޻������9�.�b` ��PW�;a�� `�ӌEX��:^:W��*�Oߑ�?`y�7f�	�WXi��u�d�<�r5��جQ���5^�{S3Pw_��!�'����qc�W!}Kx{�,1&	�$�@ <g����'�Qt`���7�����4�������5��7�sF�f_Ͼ�M�����E����Ԙ��Y;�����t��sl� ��ƔL��B�+��7A�!1�-A�P����O����i�������/��U�ջT�8��f�Db��>iYTK6�7�!�����>�s��� ����J\�v�Jk��{'I�\�s��~:�m�����y7�5�~�@����}�1`���<4%�~B�	$�7���q`��b;� a���5S���3;�o���{�� �4*K"�둤pn%\���v�.[:�l��۩�!��Lʦ�����!�x���T��i�ݵkD�B~M%Mڽ���?MD���T6�#���+��&��?�4`5'L���/(@��q	����+�gd&:c����9�C��=��^SH��l���[�Ҵp��������c�gɪj�j�V	�����]l�׃�CSU�ϻ`�$��18w{AĢ���"@͊���h�#�o�8T/��霼�`n����;i�(�O��d�*��V���en��x[<��nb��M�^��AS��v|5��g���5�S%��_#���b���3�w��'cS惙��m�2�-��q5���>g8�Q��*}�u��R��	<r�wV7�T}25j��|te�7ѱa{ĵ�נGwn{��f�g���:�O^r�f��R��[�ϩ`%Լ�ej�=�B��f���u��,�l��砞%Ɣ�ٮ|�_�8%������vv�V]iŝ9��"�e�7c&��h�Vw�\U���I$�U�ZVݘT��N"�D�VM���S��"Ј1N�Ш�4���[ �3��(_�y���{!P�����X�fv�N���~�|H�u��$<6y,ʷ�V�˽<�UW��Jh,e(�g�,d�D賠�\���X��(��	��M͚������"|��C���]��ȷ�$>�H��WAW<��C�ב�� ̓� "Zċ��	��u�ff�W�f
W� ��6��$=���+��;XD)���+��
�!4�;!�_1	t>�O<J���M1�+����m��!}�2v�K|lrȏ�8E��$������)X����X:�Y��p�Sx��tbp����U�oU���TTƙ���5�0�|���k{dv���[6�c�tTz9�����W= �Gz�@�I��V��3x���)|���ޜ���3��Y)�'�,�՟�d���2��Wa%�8u�A�|�Bٴ�v��ӛ���q�H���܅�����.!�l4��/p��O��⚞	��2�w^�N�����苷1��ÆN�(<����|�ߓ"�I�^JC��[^�E�n:8&..����Y�<�⹳�Mv�N���^���fV��^����Y��:�&���M�)ݥ�u\�Tr~=��L��.S�q�bK۰�p5��[��۫F�B�e1y�r83/q2q��/ф�3��jɒ�r�r�oY�"~�^��]�/�e�q�L�?Z�����4�+�+=��,��r椅��%�#=-8��t��	��ی�.�O՟@ު�f�'�c�J���5U��tR���2���N����:D_IS�! r�B�'؝m#���`/.�[�M~�ߥ��V�̬_R	6��5�\���F�,8� hJ�i�L0b������88�7Ρ��7���/~P���s�Xb	���U����Zn�:M
�#/Y}�[���&���Oz�`5D���n�Cp.n�0�6k�,��#%k8��>�v@�hG��ĬG����� آ�;q	Cs�����_ӝZ�@�aWYP�b.ZOVt�$����g�;��D��9��5��}�z �Ț�0�I�Sp�W`
v��jP!��.��i,��	��rc�� �t�Ek;й3�,�YA���/� �M�n?�������<�.����@���ۑ���_IF�;�}V�����M��*�v��=�� ���f�"1���;� [\?�y���g�Eq��W�r�e� �d�y��>2����1,�w�q�f�P�2�����A���缓�2��w)n�T��aw�ʝ���:VqQ�#�Nh�
��+��v:$>,�:z���o�t�[u���b�_5�n��!�va�&g����`��d��{�jEWd?�?�EI0~��N�ճ�1!�2G�2Y\���-׼��f�XշO��>[@ٰD�3`���qF0̳,Yy�*Ϧd�X�a��n�W��;�#C=�Jy ]��4���Q	�P��{�c��J�1�x-�I����d5B�Fa��R>zd�-W�Ig�n�C(�Oc&2:;���@��v�..��j8r*�xL팅̬����u\Nx ���L�C//x�7��]hRXl���w��/꣮�̑����G�V�����h�嬨�J��\���#}r68�ݛWڇ�+&�SQ.�6�LRGٺ����oY�yu�౞�+�����У5�S�V��Ɇ�u���k/�K��m�V�mS��h�bVx'b-%��Qczc��@�@�T�i<	C_E��s�>7ذ�h�u��&�k���\ �ωۡ3��h����.��v�'F�u����SRzc0�=)�r�g�<_h8egg�4��z���fL��HRcE�p�b7LqS6#�z����,<�b6���S��K��.�Bbz�H%2��_q�4�e�{|2�~�kī�̙��7�zZϿu�J�}�h"cے�T_��S����t�U�֖��u�Vk��?c��˃w������z�I�i��$V+���Qr�wN�A�����FF���+&aMӲ�*�r���!� ���[��0�"DM���^8�2��� 8��}�h�(R�*д��4�P�	\��YZL�W��|b��}6H�����om8䓀ĺV�d���ƃP������&xx�rٻI
3w��(f����$jntUپ5kAض�׫�O
A��I<���n(bT�ǀ&Y�X{I��;��+.�^�w�D�Ȍ���4�:��t�n�5�׾�p�#�gWY��Gc#�Q���B�/�C5Э��Mp�����z8�9����D�&��Y̻�����鑦ڔ�s�-�0{qch��cam	��TBX!J#�D*T���yU#���yĤ�`��.'�����w�\,+�#d�_��q��H�ǜpg������y�����w���|��������V����X.��v*~�R8?]*%cx�
�'���w�׀s�g':g��q��%���l�h��*�
��5�a�M�k�!���v>���ˑH��*���~��,�X}TM��$?���÷^��^��Z��t\r�'��dt����aӟ�?�P�!��EED�jRe݀~���q80����������G�Mʝ�!���Wp���ŉQ;@l��-~�ǖ}���5�	�ɗ�%8
�w\l��iN��S��œ�Ls�g}�Yx��]u"���k����F��K(����Wh������k j���"�U�`t���e4�x~��߅�m5�f"���_��m�q�MF}�d�o8Ф��)' P�@�/�
$�H%�Em�b�Έ�w��cUyГa�n�.A�>aUlu���.�v~K��[�*��ܐ7������ā��Q�	�{���${}���Ǒ��s�֍okk�=�[B�]�ƻS,���Vz��Ws��e��4��W�:M���(�8z��p��'�?�Ql�����8�:��u��ĸţ�,T�i��@ �դ����Aj��&��@2l�VI�EX����Rk��P�3�x�O���_�@����%R��G���e,-�͠���-�W�������!��^��1K)�}�ޜf[В�8+��������T��a�r��[����Z�W�s�X�Z�n]�0C?��wEh�����2Dp���}�Z?
��5C@������Ȑ�e@yQ��q�������q/���a�L�ұ��a�L��n7���cLʅe��ˎANԵg��x[ӭ.Ou��+8���\��@�W�2����y�r���`$��\_%�y�j��:U�^<�w��o?}��Q�L>�T.]<W�6i��n9�)ߘa�
�M �o���W�3�/=%�)he��A�U_( �1�3�V�i/�aI���ۤ�;>�	'�0�����{?��5J�VNa�jo�C���-���[G��RX ����u��=�����p��4Hj�¬��V����2����[�๷Iԩԁ��4l���bU���w5 �&ۮ�+���V4������N�6��מW�N:0��_&�E���5�˞�1����H�����X�\��c�F�,��Q�����ʀ��]K��DeU�<*d3ޚ�z�_�r��y��E���3�6��ș�� �����N/#�]kOӽ��9��I�S�wcA���Ռ�L���5��J�J"-*F���6�:�1�/y�1����/������!5�<KR� {���/=gM�m�\pӚc)+��w���8�ςe	Pj*���BJ~�谮0���[;�L���T����V�!������:�*V��C�~�V�Cy�S�Z
>�m���_	�?N=yT^`�0��C{<!9&�ժ�i�B52F���l����4脋�hgl�� ���[�
�1�q@��D�Z�@$�����	 ������6j��tp�1��)�[U���TR_����peK7��d�tU�	�jtA�F�,�^���3+,���	��G��9�tr��nm;h��#6��z~�xU}b��8EVi�~�2�g�3�B����i�����L~(cm=_:P�C�������\�`�|�y�*��z��2Ƕ�>�����#�	HWu��m�j壦���4�G�d���N����x ����fd�l�A���*��)�QԠXE�c����i��p�S�Ф�}���7�v8��^�{U��wb����w���U���l��Z�U���>��
�ô#���u5�!��\����^*��u�Δ�o�d�쌵aJ��̋��O���U5��X ��4� P�:����=P�����-�7C^(�W\�6�}�s�40ے2�Ƴ�6�6��g�4�!Y�4�m�%�PE�o
�"C��Ah���\�Y�K�nO�^�Q�}N��"\��C^&E܌�`�;@?���z,�X�v���vB�$��lε��4��G�s�v�#!C�����6&�x�ϡ���(��r�Բw0�K P���)Z���#�.����q�
Z�3m��n����5�N��Sr��̴�K�<����&�]�o�[&	�0 ��o����Ь��{t�ؓ�ѠL�D�*W���ۆ��p�g���N�<�3{���J�K�ǉFvHd��\�1Q����|^�;�9VW�DY����G�4c^ޱ���X����չ�/D�*���nH��_GͬZa�0�����p����d�AtJ��lH�^E�R�^̌�J  ����G($�η�}�`��I�`�;�</K�s��j�ϯ�c��x�1����,!��}069|˥�M�y�(e�H3Q,��LC����yb5�Ur�H�m��U��o�jSD�Ck����!Q��x!�T|o�ޕъ*e�Z�/t�Ĳ�k��&A���O�nvmO�=�(R�#p��/ZZ��.V=�٠H�c���d=���_�ͮ͵��ドg�N(��V�����*~$�ݢX��V+���[����Q�T}R���T��h�Q�MW9���з�r��nh;*I﮴P�v}�-�q��{}er4[���bU[=��Z)P1�7�㚢�j��� ��M�+n�M{ ]$t����j?Tl����
�4a������)y�$��֧�������{�X�;��Am�n��@�jO����[�R�P��'�O�� ���&�o��}�����&p��!	�C7�K[۰�~0�XYW2@�2����S�r
~u��![è����®2��%�4�t+[�J���-ƀ����=�����f���s��ǖ��Drw��O�⊫���Y�,���	�*%Sj��iuMꋧhS\!�"�%m�i�Z�ܺ}��(�f�w���{��,<�;S���,]�Y#�D�c�R]V�7��Ol��������s��>;Ż�hZEXZ#��f�=���ΥI�cEΙ���*�j���+'��yS�_�����	$��bZݷ�`f�K/ÃiM�R���$����*�YN{Gon���E>Nk�_n�L�N�	��� }���b��?����e�J��Ne ������u�>����Kk���k|�� *�s:��h�J�[�|��A'>�7?£�s�=�b��	�\O�����` 0���+���As(�BV >�`4��ߠ7j�6yv:�҂]��������p�u��9%��=�qaԡ�X�K�kG'W7�Yj�VJ[9��C ��e\�쑥߫�?����E��Yn�j������X��,�G\Vv��,��`��Nh|�+,8��'���Zu3��]��s�l����<U��'�w��U�U_�0pߠ
���x&�
!ᄓhU;؜��E6�R�S���O��d�<O�:��_BY���n{����;�{R��?h�^$�.���ew�X0��Kŵ9 a���'�/��P\{�5X�3��SWT�}d-Om^&Zbh�@�7'+=��$�<�����6#�`NI�A�鞟 %˞`��@E�H�΄�p�W�E�Z�[��~��T�}�84-.���7_&Wd��ɱAd%���!��82�?+����Y��&���_~� �m�H͛�v�/��+������UQ�e'����n�HNqF�8%{.��&uT��1��b�IP���,+����P蓒�W���뙜�t�y���*�4E|esq;7�2��+R��]����D�H�K��o ]���I"�����[��̣�[��Rپ������X�;�l���k��p0#v	/t����*�I!��C�Y֊� ǟ����L�Q3��aUA�L�9�C�����e_��C �j�1�T�}d�u�Z�.����:S6a�ZpG���G6�C	�R���U��?_��l�%·�x����H���ć��+"�� Ӽ�O\�\U�}9����I�z�!�5Qg�o���f`4G$"Pu�����"��)W�s�#ϴ���B�zO�Gr���m�)�׀CXuL�:��qX��j{^�E!����Q�t!God޽v먺	������� a�e����V����%yL��I5�B�?��-��7�w1��R�����-��u�m�0���W�Bd�"��݂�j�)� �k2��K�]J�w��B}D� �����M��(W�h��|HW'��"e�85d�(�X���d!���{1}�sWR�ų��ط��9'��`�?8.��d=�ے��7��1|+Ŵ�B<��l��>����ximo��Y5
�]���e�f��%r�>����H1�̓q���=;e-�&���{x��t��#�����e�"�8�����zk�Fx�v��32� ���o���J&�g�"�*1�e� b(�'�Ƥ<�����W_���=C����]��y�a#�g툘�_��d��~tiɳW���o�.��Qlj���b�}�
)���z3��Ovp�8��8^�lg��U� ��T&qa(s�v���4��=X���k��Jΐ�(�re5�4�Q����Z��cSY����(�c�y���ߊ	%� ��͓��궧��#����Y��H	�S��U�͓���`�
�qj�}�Un��jQ���~3��e��g�7q4e���n��`@�`ihr�g�e?���@W��,��8����ao����}��8B�����o�s�cY
��$Ӡ��q��I��$S�w�Y�8�:�}�A�@R��R��#**&?\�ʸY�u��0��� �f����1��DRi_[���s����f7�������z�D̡���L�d��	MV�Հ�	�C�o�W�bN�ڽ��cAH�i���m�l��tÁ�����d��B{%��'t���(T����WZ����jl�	��j�8s<�h�&xx�"����`�-�#6��IU��w���*EǍ�Sj�b'މ	�O���(UK�"������=23��!��@����4�j�`[�^c���U�O��/��4�P�BJ;r�Eu�~� ­uGC�y����pF`�9̿�{�+�����t�8KQi���g���i,���P�x4��Chhz�X*`�[�`���S�>�
e7��P�T6B�J����qD�gB��j��#��$t��41��ɗ�
�^V�Qm�H�+IY����`J�}Ė�v�%��z�6��P�)¹�@,{R
[�s|�Q]+J��f�rWc�_V;�<U�BJ[K�ѽ+Ơ1E1�Ƿ�"�"��%-�u�4�'�w�K���.^E���H�X���8S� �m�� �����X�h W�w��
s�C����u7V`j�u<s�tA���r�여Kr&�=A
κ��/Lxd�F����-�*�L�(3]j{ �]�tѭS6�(N�Z�Xͭ�4��UΟ�?!���n��c�染[|�y���<�'rl��,g���x��z^�"4�#E*�+-yջ˂�����P���-y_"����~�R���x��F �lg�Tj��p�������<����s;tVJ�l{{��� $�dt��H�d*��DE�<�[ѫȺkt�#��:x��p�����B�[�3�>
;���r�W�c
���0�FR'�X
HD{S]���t-����n��\`�?���V#_�.UNd�O��Dބ}��A�Ym�2��m��X��w:.$k�kc���g�vY���q��?�m)r�h�)��HG��2�������Cw@�Ԟ�Kݷ9:(������.�i���3�r�P�K7�>�If���誢;f&"˯���"ɚTw��V�]�s_�b2�����w�P��FV�l�kd
�'.� ��
��� ���s5�LP?�JLպ���8w���'�B�������yP�!VD!O�|���Z���~�-�T��V%���� ��}0a��->�Ջ�Х@%�����z��}�DeA����i�sM�7|"Q������%��U7�Lu��?�X�>Ǵ�nO��Pb�0�#I-�����Df�|`���Mϧ{d �i�I+2e0�/2�G�s�6o��!�Q��{x����	oj��ȡc�(Xw[��<�s�V�&7�߶�П���K��<νZ��(��V�l�?.�Z���=����Tg��]?��б������*���[�,o�璚�N�羈�)���1����iI��WO����U�4Ca����9|���gI���y��0x|������s���iYkkP�0�R�Hk%�Ϝ/�I�N:cg�}�c���g���b�.�{�	NmU{*.OD��j���:>yA��M�+��!��`���q*$��1�js�|N�,{wFPY���#3��Vᢋ��:TI����}��m��3�&$`u`��9��V��	{�%���%�8q���.���M1��Wi��W�-�1H#�_�A����T�6��٦=7.��".\�<�Ђ����Ñ���S3��}��,R�cs���O���� ԇ�0�����$1��r�K]��`_O{q ������
#��ޜCx��M'�o�	�.�}�E�α���o��C��~�|,�k:��-X|�h�p���%�w/����t�3���*	k���J�G;�����;�4�v���/��$1�������$�P��V$�;��
��+ Z�H�$P�n�U�m��x^��'�u�.&�d
�{t����p����%~1�p��g��w��_+�\Mi��*��q��?�0���6î���.��d�����#V[4�D'w���ѽB0$�{�2���N��F6�A�('��U����{�hV<����m5��)�SÎ`�ǟɚif�	y)����~/1������ q��E����rhnD�(��ea��W�"��3�4(�{�lvGWX�ަ	�B������r\����أ�+�{��S�!�fQ��Y��F�K��,��%�@�D���=!�΢��X+���M�r��߳<p+@�)�Ⱦ V�6�m4�-9�zTN�M�^Q���V��a�$�s7K �(���P'�}�A~(8,e�����n�BU 	H�bQ�m`��$2`j0�q����V�Ͻ�)��t��k*�S]�۴��ԅ��4`� Œ��A� �H��ֲ���" �pI7������7P��vT���)_q�ĵ���p��>D�)��h�y};QX�q�v��nL��ZG�	�`FC��/�^�,&�)�Պ��+�E�Z��7�;�ze�/6���Y�e;���f��n��Ұ!uD���0��U�m�!A�-U�X*a^�g�Ŵ=r_�5�aק�ޯ�k�X�ǎ��ԫ_B���R���$��MuL,Vg$�yL'(։��f$��> eG��\Q��_��(�Ξ�6���i�mf\�Ȏ}D�六=�`p�|	�U$Zs؜qT9��q|Y���&����T�J�Z=z��e>�_j�>YF�]u�j�iw�4&�HI{�J�'��q68M��W��������i�.nٺ�q�1 <h��t��b����tч3H�Ӎ�$
7s����t��1yV7]τ���+����B�:Y;?�+�坬ޞ��\��
S�E� �,m8m�ۺ'�ն�bL�έ�]������v�g2�Ym\��?�����e@�Tc�Ų�K����'Մ^J
KH��-5oQ�4܃n0��S��n[:OkA��p�eׇ�_��\���I/���Lm����U$>����l�6Դx��*�a�Z	f��9��*�U�!C��e;X�>7�PE����Gm�ފ�5����g��BxJm�eq3ȑ\�:���A�OUvu�	DJ44����%v*��p�)-v�"L���8�}Kv�*��e�֑}�z�I�a"P�44���~C�ݏ�|��>j.���M���7��2�,	���c
�Ό�H��(��4k].׷�ߘ�&�o��-�*%����ʼ�������#��\�����\t	���S~ %)澗i	�~��j4:�^���2�8~:�Gײ�dǿ���x�J^7�Uz?N��������'�2�δ�į���,�8Q���B|�J���Y?g %d���"�0��a���'����s[6�Jѣ;��5�63���ޙ��Mp�i�̋�$s��+fgd%a�N�i���h��Щ:��,c}�<H���ziL̞�6#9�r�e�s����a3����-��
��iu�R%��ۯ���: ����#�j���>��!ݵ�E7���"�%��F��V0�'��8�6���Z_�W��DLe�^J��o�m�@�$��&zG����e.�y�������������n��L_wt�"U;f81iMSWȔ�?m�&b�_�f4��6 �ZQ��`��nJ�Bg~�����\H�b�r�|�x�����C�޷�QC��{�x}�=������N%d�0�
o�/"��*�*��0Fv&Oy@@��>#	�Pා����jr�ߌ�2Q�z΁q��~{����?R-���Q6�F������ͺ���ԙ@�R/��/�JMg��Z2l=+>��}kbL/�x��t��L�
��[���
���>ui�QP��|�d��K���Y�6fm5+yɆ�RApC���ɓ��ݰ%(;T3�#��]�j�ݦ��*���&_|��_=)���?=�sKv��p%�t۞sY�)�?�i4�Ƚ1dT���,��:�z3JDz1/�ޔ�?�A-�w��F�0}�[�~y�I���Q3;�3-U�ۡ�)�H��Aum�ֵ}�>Q6��;�U��B�^��®�Lf7��Y	ط(޲D7c����4r��qD |�Z�o��s�%\!�³�D2~S�h���x�l�\&���'��M����4^�m��5X�"V��?��?�v��n��@�b�fsiR�w��Ax�P��7D�����99Ff>���;��P�J���.���{]�V�r��rP�n�n�(h$��'n�%U�&��c��2�R�v�~�j*H��+�7��?���'���>-�`���S�qi~_�Qk@�ev�{�9j���i��6*�2I���rO卌�Y�Db��G�Z�h�/������	�8� [�0ٟoKay  �F����"�3����r��O���.�|R3�;��h�W�c����������.��b2��fsP5:�mӌ�j[
KRc�F�5��""���d�$3�$L�i�*Ь���� a��=
	�g|��q���Sn~۾e]\�^�mj]��a�8����R��p��Y��,STe�`��E]8�B�y"�T@�)�:R�t�h��!�XE��SJj��'\�ZM���2�!�绍M��Y�c��j	+���l~P�@�8���e=�鮷�/�q��/�:��O��6�0+��I�3D3v��7Vja��Jv\�c�|�	.Is=�+
j?8�g��_iMT~�����܈v���=B�4A��d/�G��pS?��j���zC�sE�Ț4:$�W�5�Wr���	�XT4v/8x���H�H塰�T\־[�.:r|�Y��t��yʟ��5�#�$�Ab�s��*}���
�\��~��[�>}�1+�8P1��1o�S������W|��DCqH�&Ӗ8�n���L�!�r:"��
�0�G,H��Nﬕ����s￵մ�ԟ�>����օ��'AVo\��$2��j����C�P6��o��B$D�f6��}_�#�F�����Ÿ��=cX����7'ZV���)�8��R���+��mc�=Bἔ��7�����g	�l����(���8�p3�L�Xu����b �粖��0_��3V@�&�`�D�*� �����u����4u�i@ysF"dQ��
�l�gPl���Vү�C���s�l
`�kX��}����`.lu��Q1*ʽ�Xy�?���΄�*�Yc���ti��ki�AX ��� c�n��?/`�	?*��lB�F�L�`ee����#��`�no���k$��0C�0
�w��XSR�,���V��<�6\�{�!|q/�����GgQ���XV����&y}��>k�Z��K�
$���ȯd���P0U�Q]��$��k��\�KH(�@��Q"��p�x�Oķ#[�2��
*�?d��LT����ke�x�Ԋ�9ϵ6Ri7��&j�a�'~�+�������H�3�D=qC���ݥ&X��|~�����@U��̋����{�a���g��#���
�}'�_��?u�N��z��ulƀT ��d�u4�sr#
`���c)�[��;��ی'����a� S�M��X?Fj���|����z�g綞eh�|��A�@�Uua����k�O�X6���)�������(@2=cղ�.9yVq0B�f� ��W颜Ěe�$ 6���#��?m2�-��!����Mҫ��d�N��p^��s�)���BL����/�Ӊ�q�����d���#y{V�Ί��k�$NQ�����Os44�hK���n��iw7��/�ϝD]"���<�_�!K�9����߬M�.��=�y��۲�q�t귁mb����k'4"���E�0��a���m�Rܶ2�X�$�ɢU�1)[v�u;7�Ē���Qɷ4�R�Yock��?@���-X�dg`�Kt4�A��?,��;Q���? ��66�W���
C���A|�okL�"�o7�|������ᘺ�YΙ>F�� ����'�\c�7C|��P@��#@E�{{�OV�e/p�X�xs��/H�r�Ǫ��jF����E ����g"��V�*��D���w���
��ia�|��!x�*��Hݩ��.�A���ӈW�%CY��$(��4��3;~�o�7���RR�g5 ���0��!���'�泵�󤎺�5mqr'�,�7����e�uԩ��kP.��hn�.�<�h4s��I�#��*�^P�( oxǐcei��:���Kͣ��֚C���0QXБ=s�W�7�����F��kR����Ë%{���>D�� }��2P��cE`�C]�R@M4
Q�M4<�왨1����
��M�e��t�����%�b�!YhC��&W����l��J����l�jS<n��V�9Y/Ƚ�� �&ר̑W7����ʐS���i����!�Hw�;d�HA�y�I���� (�\q?	
��g̢;��a�����?t�/%%l)-���m�S�r��Ux���,�g��w>���$��!zvXA�Rҫʮ�	��p5�����!co&��*�`-ڥ��7 ��4 ޥ0�A�pH��� ��&�k���A�rX�с創��	���I�@b���39�����bp��D[���)����O�{д�6������4�]�u�n�
��{�c�L!��C��z�_/g((�̀]���z�7@����g�F��5+��n��m�a.�����2x?��@���p9�4aZK�SFr뙴&�
D8$�t��7r�@�Ha��9m�̋`����*nT������AH�=
]�/�n��H��	�vԍ�LkC���\>�xQov�g\��'�q��،A@h�^��7,Է���)Иk����b�u����_J�UD�o{q���`�g�!��d�� `��j�(e�;�c&�9h`
5�-��qrD���uȱ,ϭ
'N���#L2[$��KO1���_�*	�l���!�p�!�[8�Z��!�E�š�e8Q��7��
I��k���K�5$�]��gэq����Oɷ�����_Y/<��3��������`�w��l��j�5�2���
\G0��(����m�����[�=0���û�9�������Z���˦�N��d	�K��o���8IVK`t�K:��6��1@	!���v[��c~�RnKc��2�?(��~���v�b�a������0�)��`�:W5O���㫠��ެ�e����2�N��@�Y���E√��Lq�WM��>�
���mj�����\]{Xa/�P��nϻ����l���Nb2e�_¸��ek�_�껃��q[2P��0N��V��입⏸gd58�ȘA�.�PCNj�W'Q�E�@(�[����DY.(P�1g��\�����_GL�l���w�a������~P��[O���ngceĦF����X��:,8�������ӗ��SJ&��x&�ܭ�i��8��Ac0 K$�����	������R�w&�B76��aMx?|�:H�����A�[8����y���~<�s���lO*uoB����vK��Һrd�|C��#@�'A	����h"��G����XwNʫ���L�r�H��/2T�=u�n �1 �� �î!�NR��E������FG�1ⲻWKD0^rɆ?��F��{G���e�߱pnl��Ѯ�x�-���)�.���W�W�����o[T�^����g� zf:�x�]q�:\y7A�5Ѭ�BnvrU�5Wyۗv����t 󳬹�u�6�Ԟ�[�R�DpVM��:������/�s�X�yE�J�}�rC0�S�Ɇ9z���K��~�Cݚ�98�;�^,�-��K����A^�i�N,":�yJ�е4'"��d��XWN4��� =���T��L�`cka�៏g\��&��V�k�Z��ƻ	k��G�Xa��ʾ �e�u���P���F��Kh�GiG5ަq*rҨvvy�89 Ƿ󔬈�6gQ�_m(�"T`�����G����/�p ���\�6u�̧ƴ�_`oE�:���%5�=6��C��FTN��ts]��Wݔ�-tH8�NNr.�q��(�
�g�S���+�v�z�3����u w����\����@��,(���V�����UO,�ߚy���6<=�!�6B��x��{II�'��t��o��h�qŖKU��5%lY�۠�d��!kg<Z�_E����x�O���a'�����4��k�9ʼ��k1>����е�:i�z"D�#�ȃA���e��n�2C�*4���H��
�sOJhb��n��}����0@ǯ�˓�!{����4p�uV9e�Q`~%��G�&�O��t��[=r�b
�zt�̋x0N�F��6}��[e&��u�I<Շ�4>�WCZ4�yzFq��m��D�7m�f	5`�&%q|���,'*J�ʇ���2�E�
���B�aSο�~�����Rr_�/=a��w��r�9�j�Є��dR�C07���"8q�!��<��0F5Mm?20maa�g��y�l�S9N2� �旅��o+lz��	�}��	 ��I푥��J�-
�|W�%�.�k%t�cI��^_�g-B7�ԑ su��Fs(�$�~�#�$��Ifo��v�X��X�
�VJj��T�B `%+m!N�GW��pl���募���~�u���^f�e��ej��X�����8�iF���RR	u$�(;�ŀ�?]��.`�»2����*	�t ��.�!0��Ui�C��V�2q�Q�˅��9-�q��������v�D���c3.	�|��$��&�g��8�4fv��v\'����'$�G�C��z�D�R�L,ŀe�q+��������A�,LIs#&@f�,�w��{�ErV(�{!��,Vg�~� ��,kyYG���|�A|`�1.�����߯�#�{ӈ���TE�-:O(�Ed�-�X �U�G!=qH�Q�?��F�����$a}M�P+���8�7ZQD����s	l��"��Q!�X.妇d��e٧�<�{X~��vX��jv�֓��͓�X:�x$�Q �6����ĩxd���ͨ��'�{��%p�!]�I�iW=ހ�;aq���&i
��WK��[yQ�G !7ʑ�I�[�t�J�A��|\̩�WE4Ѷ\?p}K-�Q��'��H�A}�v0�WAs���KL.پJ8D�����:�8,k[���� '������|�[��x��q���Ku�+���}����S�=7��p߇z&�N��2ǥ�`�;�k0�
�q�ݍd[�1C;��lWh]���n� (�����%#lċ��0���*��B���,�&n��41�e��%dn����%w�04��;��\jV��BV�*��G�j�[au��<I�gowPrڿ�j��.�d�#�M9�R���2���'
��Ze�h��-�ϸ��K���@�7z�'�\Ч��*���g�f�H�����"�aq��5r4ߎa�4����{��x��n������i�`&���n����@&�A��W�u���.�-��G�Hұ.��#S��;£�̜�(IOM�T��q� ��i�6![4B�?��A��_07�:3��m@��m� �[`m,���E��:�(�3������jJ5���@ˁ��_���3�N[Rl���A����9�OR�\N����� >u%{y.����^��/�Pe�t]���{��fފ0��Q ����+��6���Tь��@�%w��b��X��丹�@�ێ���âT��>�!�;��ҧBϚ2����3"Vs��p�Nl�Å������M@��q��G<�k�t�������@T���`����.�잢�����4����J�����Ք5�q@'�8�$�#�5-�{��>!�o���SZ�)NJ0w�m��|�-�ۆ�t����P9�e�\�,f�?r��`�dL��	�e��!7��"�.-*Г�Ʉ�q�Z�m�����ou@3�D�
O#��lKwh$�,?R'g�G"��^Q	d7��/g4n=�Z�́?��ش�_y�Q)����ڮ���L�N1 #M�b�$
r!�{Ƒ^Ǩ.  ���xp}������,Q�(
d��Q��99�N����KhU�;�f%�Wxj�@���k��w3���� �yt����t04��ǿ�<�����5R�.�HV�뱂bA�I�(���;	�U�T|?���.�@�VcȤ����&ƙbH�uS�'ߍW�j?����l�)Æ�Oqv�d�����뺞���6~�=��w�6؛���L�?}Ϧ�YP %@;�a�A���-�YEmq���$�'���w�{��Hl�V�]
�w�����[����M���rw��:( b�|�S���}�x��#�������Ż��I�(:3���JNN�D��jC<=��C1���0uhz܄�TlQ��V�S�0�]�_r�>B �EEQ�Jz��*^w<��RK�ż\��?�iC*Ϋ38ֽo�n^�w�`�_��q`q7	s(b�\!�^T���Wċ!_X�����!ב�L����]>'�uT7\겪�!?j��M|��In����nc�<�ߤ�8�~MDVd*�/*��n�~�pp�����o������n��D���
à�k����"��2�afOG��Ί���$�Dr��iB�HE���1Dq���?Y��(���^���a�2.²�=k���ֈ�n=��q;h�jcDe�-x���?��j�6��k��7������>�[���>;�g�ٲ��%T�E�AT��$JV�Ӫ9���,��spy~���R��*^����L�&�-��]��C����U��J�il0��
k�b::�G�k�}�	�h�:�yT�z�疇�����3�0�Q�NX�ZL
G9]��u�@ڴPt`^��'׽8�"�ř���Z�ҝ+܍ju�)���W �(C���*Z˝\^,ϊ\f��V�Fa�r�K��6i�ֿ�t�Z�L?x �[~��{[�wf9{��5(H�2-\��c�'Z)V�pdڛ�)OP��ߍ��Ý��޵{��h��u�������T�߮�$�'�krM���P�b1�iyV����:��&MS��p����lh)�����W����C�L�I��I���ȥ�����h-� ,չB�iKs�E�)��p��{T�狪$���^�fr����8w�w�&jn�v�Y(kG Z���yrW����������4[^����� ����?g;�f�|[Di>ʸ�����)�{Xy+Q[�[U]23/=-w2�rBvޖ�1x�kZWo�&P��Q�����3��	K�q�2��J����?�B3��D�'Nw�r�QE
�å8�vp����+�MKZO�	����LrQB��ԅY9���GK �˻��X{��=�"�n�"�V��ט������D
R��,.%=���\�V��̈ ��m�o�^��� �f<�]2h�U�.�����$���u�m����]����Ϲ��/���1�(/�n�W��jw5[�"h�؊,����V���&�����麧��d3��.pȄ;Yf:��?�%�C+fT=K4֑�V�8W��䫴�'���r�@�}
��% ?���,Ӄ��a����_'g�� ^U�+�Uq]��z������@ݥ�)P������@�K�5���R�S��#'o����v<�]8.Bb�4k#!�g+�Q>|5_�OF��~��q�.����,��z~z*�0:c��v�HU��c��-�
��,н�}����a_�4X�����"�O����N�֨ۍ��^�]�������{����4ۅ���M첊�(�bMu�a"G�;��|�ga��t��%�4�3�����eĥ0�a4�n�,�q��%�돚6O��4Yq0f��Nc��0�%�-�il__WL�A��'�^�6X��@~@�����I�2�ʱx-�kY3�=��#��������,��$���W��	T�vt��%a�.)pML�Gݼ�y�<�����ܱ>j
�h1��m��ዣ��y�C��]&�j�2�gOH�;��g5�7fW;�85���gӮ���J�2_��r<S+����|�E)#ݧ�����v�ڳZ�-�6?p��������{[��_�ש�/+�@Um�3���4%Ki��ðo�_	/cn*����U����u�Ǩw�J�W
�ۭ-����{��� �K)!�T_m(�
X�ŖȘf���u\m4��&��u��2bk
�ʧw�7��K�7��r}�֌��:�����
`�OEP�4o�\l����j�B���g���|�^E�ɏq�a�U�ٝ�'�X9���8�"w0���T`g��Y"@��?ۭ��ᓼ܅�K�V;՗�J��Ί������5� �S'l���O[���W����"v0+KB�PBN�~*���̓m�@���iYVG=��BN����r��X�������\���P�˾k1�_|!"����-�����T�o� p�S����r���
�צԻ�#:Ф?�-����#�18�\�k��L_!�`l��W�s�eY���'�bJ"����B�zۜ��j�1[�?;P�h }���'���!�J01�1/���uU�����C��XR�׭gzB+���l�̘�^�'R���m�7��{a$I�þ'��L4�6r�����v!C�b������k��_#���X����Ÿ�5b&�x� �~ڑ�		�Q�L+A�(8���4��Z� ��0��{�{C<Y����x��;L$�V�]ͭ��8w��H�U�X-��C��a{�3��t��h��x���v� U�l�
�E��|�i*M��ή��z1�~���e"ڵ:r���Q\��{�.Y�CO����\&�%a>���E����+���73 >0����@;�A��I�'`(#3V0�ō�6����=T���6�]���m�^��������c�65����y(!��҆�_��t��$��uKm�?��=��\\�Km�OiCK�{�zA��և�C�2�Jj�6�N�~��g��%���[ �F�쩁$���nU7d�	5������:p���t����̌9&p�OwV���T�aS�ݜ�I�d�V��'q�[C���s�AX���� �`?5��G�z�5�Zo�6���VQ^B��ĮV5n�ȻK7ʯ>��i�f�pY�g�v
��
����Y��v�0rh�QE\�8�h�8?|8�U�\�F���dn�t;��?<���5Ԭ�
�k��o$;ߎ�&ňV坮c��BD�#G5���wxj�5��ߞT�p�n�l����������ci�͚l.ސ�$���P>4���Bw�m�̰y|mK���/�k9
U�O�{���]������m���#������^���)��Kղ�q�I�_� �^�;��zJ�W�9�dE�Q�g���޺H���f�7��*Y0��V�*7�8@���)�yB����SUɺ���@z�@���V�<?&4i����B�X�ܴRs��U�� �R��gwǦ���i�'�T�A�L�u��U�qf
l��Ef�(�*�n��*qQ��r!����;�%���Ĳ�5���W� KB�D�]�����Nl�UsTS�-C�N'`~��p4jK �hѱ@Ko���T}t�Gԯ�$�1n=�X[)b�r���$���*GZ�yD�>=;�����H�>g2V>$�p($P�㥔N�&���_�[�}$��<R积	$��'Xa���t81İu~�Y�2<��H����׫?��shh/
_���ڸu�(���j��J�jN[���m�E�L���<��ii	�9��>���Z@�r��%J�j������7��4\�߾���z���1����G:�6�Q�m�x��I#�YE�\qW������N5N��.�[V*��M��Tiy1������7�����+�#�VF��%�M��#.H�hk�Bj���t�ʴX)~w�EUR��#�a��d��*!˪�(��&�CE�<+��ٛ��>'<Ğ�
���H�+�\�9�}��j��?�q�[�
_ �~ ���M{�{ӇuG_�̣/��B�����]�.�9u���qgB��ӫ����I����_�߆���H��- ���<� ި_��ݽ����@����c������6]��P_�L�<��ix��V��'�7�k9sV �5�cM�k�5Gl�p|ʏ]��K�2��`ߊ��b�ԥ�=���-��2��e��¶��S���)Rey3�XC5�J��1Ezha����_h�v��a���YB�	��V���jԦ�'�UrÔM�_B11v�f���ˍ����
z xOpn���M�p����@�H/H�?z�o��ұ���Ia�Ew��G�ʙ��]�cG\���_{lV�����ev3'M+m�ש��P��!���1P�K�p�³�������ܞ B )OP�أ�-��I	�������k��|仴t}��G��m����LO^\�1������QEC�d�\_=w#+�Ƥ0�K?l罸@n�w�u��b@#���E�J�Gݟ�~}�z%�����d¤*u	$�Ǿ5��kB�U��3'�6���$X�f��-Gr?�$V�uV`~���(,��~��_�C��\�S�OM�ߣu5C-7�dR93V�	��b�y��^A��).b~�.O�ͼ���0���\��z���˵A3���P�p�B�n����Z�m{���B���mz�/��p�������v�N����"#( 8=������{8 ��V�o�s�KXI�3��rUE����/h��1�s��n�3g:iT5���,C��o�� �$�|Ak��va�B
�D�h�9P��ٵ���N�P�4=�/��Q�ui������~W��(5�Q���2�?���z�f��%�8�����j�(��_1����N������T�=��}qPJ쾷2��Em
^OM���c�P~�sv��(G���=e�Oq�	!N�����V��������GG.�������/��������6��G�e�r�'���[�CV�� ��hvZUs(c��?��[/�Z4N.�FŧN��$����+�����-��8.�	:������f��\[��-��F[����}^�!�CZ>���Y�aH����K�I�:Nㄨ?^�"d=K�Vh��ug1����t�Q���1���)͛`GF��L-7N��@�Bx�CyEw1�K�jLD].�q_eGM�	�o����Q+�h+�7~�:q ~�@8H��'B�����~��;�
`<���9D�9_��"�C�?��m���ь��ѩ=*�Ʈ��B��a`��IhQa[
Qa���t���	�C��~��^��Vԩg`�����}t����mKp�E�pA�5���(���X�Ȋ'g6?� ��r�4Jp�u�����aю:n�oD>���\�Õ��8��R�汵b%j����oO�Z�[3�[�p�i�s^�#3���ؒC;��@�8E�,�^��^���(�D�s�/|��0X�@=���׻/�Z2�CkR.qnW 08�J\�:C_pf6�'��J]�i��C�o?]��G^b�u�1xd���'��Y�M�����?S��z��ݿ�z�p���G"�)�_F{�L�s΢AIU�U�� �v��Z���$G����3eB�o��˾��g�x�π"թ-k;7<�����Hq�kOqX��u��԰=�- 9��=�$_�ÄL{fZ�|��'���jS��h!Bp������˯L����B�}xg���}�4;��c^X;�ʠ�>y�u�.8׬SI?1�r�JM���r��N�=�����;��C$����H��h�wT�m=N��Z�B#n�`dZ6��a�2ͧaF�������[S�\�����z?2�k�A��p��1w��6�ul�&���(-�2�
Q�b���C�9F�=�fd;Jh��0B��>W؉���M��j�8f��O�C�e��� !ܗ/ዱ��������o��X�z���H���P���r8X։�ݤ�)1䢠�7Fg~a��[�]j��+ ǈ$��д�������T$z�p���-Vc*�]3��6<�/�w#��D��L\�eٓ:����W �@+��r!�#�2�:�����<��6U�-	&��^�e�J����sZ���X���t�C�C�4G�Q�:�A�J����un�����G����9�(�?e��\��A����ĘQ"���$�=,Kޚ'A��ûH���N��#�݅��K}5�3�$!%a^�Z<X�fsx�X�U�6��R��ſ��F�#�1����w���1<U�L_7U\�Zj�r�ǡt3`I,��[��y�%V!M���uk���䮋��@>����VtsN���&�������hq�`'��Y��Yg�w�-���~���ɗ�q��!�&�����^�������9PW,��+�B�,z#d�^tȲa�|��{�W�:x�
g�|�	��9�ަI[�m=�G�0 �M�g`�7�J �=���J6�hO��~j�C�eO1��N.X�SL"%��o~�=�K��q7�Y�P���xt@{S@[ǘ�m>٤�����'��ejbl	}��m;G�����]g��R�?W���t�`ɐϰ)9�p��G�j�TI7�&�d�p���=�,x�q��_	of?[T�fq�4�N
WA��T͊�b7��5`�����%%O<�bl��΀"���>)=S�N����LD{X��V ��zE�����7;t�0�9��i��;�WG,y dB]l���'A��� �#��SD8*�InqQ>����������{.�=�W�4{6c�����Yy�jS cV����NP�0>B����Py��G��	nח���n�o>�Ӱ�w����8�Х�Rt��j�{�/�6@ឩT��4jqYeXeX�����W��\v�x	�t#�p��c;ʴ��4�W4@FPhd ��:�뽚L��.�R���Mb�4�t)$G�b������>;[���Ȑ�'u�T��wTs?��k-е�6�h�� ���k3HYn�'�C{<5���r�]?�:��f�l���e�I�w|�6�IC��gm��+���R�F$�~���u���K�:�VR����}2V����|�z�x�n��yƳ� ���pў��c�>��J_�������B!��bc:�u�-~�Ɛ��*�>�I�U�N����$Gz������*����������IL���#�i�k7  �hفtiғwCk'��y�Z1�XKE�t[�"�s�Z�6�Oq%�T��!��]x�#��8��!�LTP%HiH�ƛ�߭�>�|��*�$[�s�ЮK�&��q������BoMA0�*G	�#��˸0�%��+�+�aQ=���S{��*vf!�@�PHtd��0�3z��NR���5��( D������0�aJ�aշD9��|�@Y,tmA��wW�TR%����ZZ9t���_���ɀ92xl�� 6�g�hF`}�Uv����h[]�P	$In�pR����VmC*����z��j��e8z��yӂF���m�,;/k��ܮl��0\V ���w�{˰Uŭ6Y��`�Z���~(X�/{'���$���Zu��$,;�^"&Zדg<�lzkcο��AT��Mǯ�-�O#Cd�Z�C��	ÃUh���A���R��;��X�*���ԔR�%�&�uD�1k���G����\��lQy�qA�z�5��k�BR/G�����E#{kyW	���3��"Q'��e�LvFP��VYw�$��	!�	ز�g����.����=8x�eE����$+�����b�����r�J�#��:	I,� b�
�c�~t|_bϻ=P��g޹�Z��>�RݏO���>{K�#�JH�%;������[��e*�ǲc��0�j�U�md���Y9�Oe��Ȫ�@Y��^��Ĝ ,������tb�U��y��,r�"��	��*b7�����=�"E��P`�s��3mt%�Yl#�A������WԞ�!���^�p �A#..�v��&cC�{��h���Ev���ۡA�<�U㸂6�nk�4��D8�\�+�t���~���А#����c��g#\p8�%g.��a�Ț�>��ZO�EY�i��S'�E;���x��v��	�O@*�������q�kN�^��d����~��	��I*P��k��Ѻ&j�i�(�A�I��80��CT.���D&�n����4/I|��#�﹋1��BЪ�"@E�s��z�.f�7�T���P�ζhy�\��+���Ð���'ܯ�['��vP��V�w�}���`��W>k����_D��k8���ױ���-�4"��k�$�Y�� Y�x+�+,<"�{˧�6�8}@�o�q��S�;Hgv
O��ue�S6L�{���L|�����^e�����u��|���ۅ��i �����-�UQ�d�\��������8����"H���,S�к��S�Y�N�w��S�.��ʐ�J���%�_Z����#.�#�d������}�_eܤ6�˵�5R�ؑ��)�6n�ӷǂ��OV �D�	Ϗ�Y�*��
;����y��֯�,�}$���E��,ӆv��^-iZ���&�E�x�aX�Q�J�"#F4�	Z�C���δ{'��>.�ts]#�hT灇����pP1�im*zQ����Y�@߸{���ئm游|I�%K���C���a1�� z����}@Lw5���p`G6�v�K?ch����P��W���Xo~�拙H��N�M�b�P�μG�td�ij�D�����bE_t��+k�b�cm۱��s����4�^A� �5l����3�i���a�*;�QCX���D́
�JF����0�?�;I1oU9b����2��ޥ���Gw(�dX�Aja�R��Q]RR_��b��	}T��"!�38c�ٸ�t,��8b�'%N���Yƾ��S�m���x�F3MY�8�{��bmк ��9EZ��,t��#o�Q��Z�("{�p(��!M�:�	�d�yR\<�SТ>��=����v��#�Q��,���t�b�1i����	������W�qrX���[�қJ�=(a��w����1)O�,��-08�y,-���a~=�^���e�Nwv
�%��YR��,[A2ؼ:��lai���Ë�ZM��g���A�����@i�'�a`ǽ���X�y���3��}�f��d��-|�ٛ�L -s����:��s
�>�c�I�A�>`%/0�e���D�Ƈ��<����@��[��pB�g�M�i!�k�ĉ�[��!�1�y�T^ڍ'�u�1p�.X������t�V&�V,�9� �yur80`�,�3������;ۋ#���a��Ӊ�W'��$�Y��a'ni�e ���Է�߷y��NTk�g�>��ۆ��+�¸,���6��,/9�~�����~�#$����B�d�>��HQG5�p:ڿ ����yL)��]���ak�{>��6*c��V�6@<��h�Yg�r	(�N�C^�fqxk��^>���BȭCE���]ṿ	|6�L���o���R x�� �b B��]d�xÊ�,��C!6��m�+���ݛ�j_yg�O�;�./��I�����A���~�;Nkg��^tD#M}!ZG�����Ԍb	��c��$�uR;�&�
/����ޞ�+Ee÷Q3�(�$��S�s����h�󎗂��%,S�U��\���x޶��	�֕������R�U�c�k>�c}s���]j���C��{�~N���t-!�8���m��?�=�\P$F>��j��rEu���>[���I�}���y��N����XRp��'$`u�<P�Bw� ��[�l %W�^=�������`��a]�M����M���Z�Z �e�p�w� �U{���RK��瑏؏9�\���Ci:�V��{�ozf�g��*�*���훀�v�%J���*dƈ��>��0h;L@�ƅ�R߬!f|���=zV��3��4�L��A%���)�H��@Ygm��(��o}�p筡�W�ќ�L���U��V��*l�bJyઅ2�tF��hLe�`�u��ŏh� �}�@���{�j����][g|�Z�Ч4��v7���v��rHH7�tað�5��YPЧ�lq�i`�W.�P��B^�1zer�C�4�90+*cA�����M�g�wc��ϳ��_�?E�"L6K�N`>0���K��V`k���42a:3X �F��p#2��l�˓\W'�sA��S��w?~*�:x�>����uH��yCj���z�[�-8EA6��}�D1\xu�W������ϑ�d Z�+_�y!v�rbn0���4�l�=:�ԐA��=G�8il�,�8�=��"yx��'o�����D2�G-��{���;4u)r�1qt.�Z��V�����o����:�r7���|m-��ss"��&u�֟�S83��˃
e�F�		f��Io�@��@�*�?���8dCZNlr⌰0�hq)<����~��V�j#�����S ��,^�#���w�/�<�l���J����!Y?��)+�N�dLޝ�W��K���s,���E� �o�ǈT�<�6�$?A�3��5����JϮ�%v��,Ǣ�������7�hk(���js�9�9/�+���,��Ƨ����Ұ��>6R_�W�N�g&�
m��a�K��߸�=tM��l�:p��A��~�!�����M#o���E`�l�WO���Vx��yA�6�6�g�7�޷ᡇ{�)H?��ܩ�����7�o���Bm�Z,�p��FC���U�W�=����J)�K��s]}��L�Ĳ㲄P�G�ͧȼ`��(���wEj��XE��:�	�qexBai�S� QFU�A���"��>�̝�����]��P�-8���Nbn�<ʠ��SIe�������޷���* � ׄ�Kf�ٙK����095�n��.�Yl��N�Ϧ���f^H���`�q���)5�r���� �5/�rV��LP߲Z5 �Z�Q�����Y3�xt*Z��_L&a'p�^�?`�zUm7�q�x��o��>��x�i>�@�=�~J������Dt_����NO���m� `u��f�ob��e��A<�~���0�ϥ �Zڣ��Z�k��6�
���	�_�?��=�F��MX�$�(� M�'�ʖ�ԖZ]k�a��Q7�N��㥁� y�"�ޚ��S�΄-Y"�CQ���g2��Y��uIdk~�Iq���L�y&�(Xf��Lt� �Xz{{��"ˮ���y��L�8y
n�U�	О��A���;��FHLu����9�ˑ��h��e��d�1�߯.��dl�^��x^d�4�jؐ�/��ڗ��B��������&gc��?e����ߧ7�V�=���m���d9zX ;k�h?�5��:�����+{�а�+�uF\�"ݱ��������Z�$	Y�鋪�`��G���5Z��O�x��$��������S�CV:�Յv�i���c�_���N�9��|1��B�ZP+Bv�����櫆C���nT	@���"ۏ���ٝ�'�U��B=RGz�Mp�z
��v�-�9���^�%&������x������2�������9�#�0���o{��0`������,���)l�%��W?��|������M�0ܢ�]���{v�n�[p���8�>n�Mx�%D����8�'�t)�oʵh|9��s/G���{nߐ�Ej�~�`�ě/���@#ɡmN�Bf�^{�<	l� �iz���m�����#B�1�o��m�+C�"~�Bn-6H���>������s�cr�F��q��W�rt7�Te�`8b���n���l�e�wݍ�EC�P�t�3�Z R�>:�g��/�mV�B�:F�5|1����;����R�"��m_b�̪͛/�~����~�-dq�*��b1��u��jXR�ϰ_n\�jC��-���烙��g�M�ma����f�ܡY�z	j�T����b��~ӄZ�v�t���N;��W\j,v���mUb/{��S}=��m���x�C%���eM'U4��{��	��r�~� C�U_H�]���Vڗ��A\-�4��I�ͦ�9z���NF*[�</�E��!)rm�gl�W(�����r� zl�VWKJ�Ќ��]�l8d�\I�q�؄r�V�.�EզB�I>�d:���X�Ze"���k�)S�+�jK����'`ҡn�t4�����h+2"F[�����z����L[�Oij��";?¨z"�U��Bұ	8+<Bߑ �V�g��H��r��HP!sGГ4ia�nJ��N[��Iq���XW�cy�5�T�:]b�!\�!i�W6N,.�yd��Yٻ&����Է'��I�[�J��7p�0]��yڄ�	gU��mC�C�!�2�w�t?���w����H��
� ��n�y��u{iH,�!i�4�'6#��"�t�9^��lӛ��`��Im
�<�Sc���\_�I }���!�Ґɯګ�:+n	�{uk���x�Zn�0����âe]?)<,�i�Q�\p��J4l���d5��Nptm}�3�SM�*���Gs��t7�]��O�s��"o���j�T�T1�P3��r~��"EK O�fl�������UH�B��^�Ǻ8e���1_E�~�\��ź���Զ���
�˒����'w
�kp�%�%Y ���Q5K���򟖛�Lxhb�Ea�g��g�ic.�X0�'��r +Os[�&��y�>����E�q�)G�[1��\�?�e����ԃ����z�K_��uwL�Ar;l{�!H�>VW�7Iy�(��t�!eW������{��� �f��n��eh���0K�W�m�H��n�����OK�h��/��:��+�|he2ԡj�Mb;�_3!X�'�r�M��:N�?3]�z6 &��Ph�csri��Nx�ƞՂ&�tY�2i��T��`�YK�@�j{GwS�H�Pa�?�Dif�(]���nk���[�7���EW���G[q��Lc6g�V�7(�?e�G�oB����ѕ�6׀p5��i3O5�q��!��z�{�o�!x�;�˖�����g�
Y�&���p�ėX�J`'d��o�&7%�)+i].�3
��#g�:n�Q�n;-dn��?�����u�1�.kV��,'�sG�QP\�R�a��-�H�b�%�y`ھ<o�ʢ��ٳ��턧����,�L�[U�D0�/���ܿ�/���0۫�q�!*�\�s୻;*��?K�0�:���`yv��,d�Z�N����rЂ��H����J*e8��.f�Z���T��r˰>�`
,q	+%��3y=����lX-�Δ���ʏ��
EE�Z�:@���� i(U���q������w��G)y�^+���f$c�U�7������T�i��H@�̫�G������;�L����,�H��B%e��t�AdϾ��b�٨���N0%��T��SOQ+y�}�0���Z��)�A�N��ȏV��Oֿ�Bs���q�jl�s���X��K�����ԗ�W��_���J,���ٗ=�L����M��#���`�q6�v�:����6!��hE��z�1S�F�U�'�{�7�9d��Big�s���þV��J����<u�dxb}�j@�x���<
�m�p�W�`�;҄�e����!K��3�h��������==�CD�����.�G7E�֋O�h�����:���#�9OYT_���@���?�����H�Lw(�2m.:�7���05��ZO��\L���6@Oɨ�7qwSS�G�x�(�@�Y����?l�P�De�`�t�l���j�����Y/YGٞ��C0�p���u���di����xP2��6�,(��8�{�B<z;��cN�-��b���L�d�������ç'jXZ�B'J9@��J��l�P����1��/V~��\-�͑nl�v����4Np�S��'��ɘr.۠.-��f�����aH��qM
�a��'n�G��L�ϕ���ޢ�V�4@>JrB6�M�� �oE�}�9�R�G�1%�Ѥ(1����uy����~	�0�=`o�[���4�b�mI��.��	�:P؅�ؒ������UC�	���<?��{uh��� f�EDBLU�l���҄ƐB@��I�tH���nej���}�SY_��m��z�s��ʪ(/���Fh����K0���l�yn�Ў����%�eu�wz�}��i�8��p5U�� HƋ���J����ÿw�C���^l�'p�'�}�V� ��D� ����*g��./�A���;��-Ȋ!���>-���ɑZJzr�r�m{x��pi�Ji)]>':�*��@���=)!x5χ!5��W��m��������j�@Sʐ�+��*���O�/5� p���sz7P���s{;�x�s���L���k³�ꜰ љ]�S��l"/ӄ%R^�
[��u��^,�:�|y�>Z��᦮��Wΐ&;�w�	H�>;�}]�%5@�.����f0;��W�P�\�#J4JH>�:QZ��yy^��Mu����c��b)C��̌�������:搑�o���>��|]?��h������R��Jr%����f��^\F��o�����
h��ر�4��p����աh��B���/Lx��u�-=W/����Xlaں�6�&Pn>8Bj�ab;s0-�I���+��V�K`��\�5/�����$�Y��v�V��#VL�G���j�0S�#�%i�ali��/5����0�	1��B�����e��zI�Y�1gS���H�}��[���8'���K���� �8�W�"��&�ǂ���-K�o�}8�G��N��>^��|*�t�Z�C�L���+��q����'���0�3�Ps����gHC��tw�#���(��Ŷ��x�2ܮz��6;��T��[NY�Z�8Y���m�&o��g�H�#2&#�����	@�m}���oP���D�U�.��md�5�/�\؇kn�&C�?�d΄���X��ԀW9Ʒ}��6=���!�{+��䊺��Tc�Hx '��2��a��n�'m��].<��K���Q��'o���f1�;MQU�̏�c�	���XH[�a�|�l��T�$m�ܓ�QQ$����n�-�w��tL.$�r0�߿M��Y�)>�����z��4`Q�yߙ� :=���+� ���g�߃ȇ����QӐ~��T�o^���b��C\�C�.�u�Jt�9J�ė�B^�%��,<�q�>��j�����MkuH�KyŽm�C�Sx��� �ض�ݹ��h���_M��UM��B�
D�"z�U[3�B�S�'�^0���������G�����y����kD4J#x��i���ED?��q�ׯ2N@�R�����~8�%�� �p�M[]:N�2�Ndt����3���q�_��(�4D�sw���QoY�D$���u$c!aq� �m �Y�&����v({�^�-���
`Pg4��)�4z���:rk~@W����X�T�0 ���	k��d�rkl��}��4���}������h�-��9N'><ǔ=����x����1���	�#Ik�u3�b�!����|x�m���
�V��B��e�̩� 'e�9���/ ��aD��j���cv�W��sG�f��N�=3�"�M0���b�8=|a����C���H�K�ZG���4�"'7��p��ok�T�����eч"ż�4�T�zjV;>p��c.��yk�=|��[,|�S�/��񴵷a�IȄ�*Q,B��W��ڲ�9���ڣ-�.ߴ<i ��:!����^sBr4�!�
$ċ�����������r�q��9��� �Jx�k�z"ا6�������<���ʈ,?7�K����RTz�)@k(Z��H��D�
.i�t�����֪�����-�5f{��w���@\���ϟ�.�$�䳊�1��Y�,�� �P�w��y2�.���Nc�Cʲoc%6Z� ���^�Z)�hR�ɍ͊ݕ�V������O�J�|�kf
�X8w	\��@v=���Yh ��j^z?徨;���Hx��ooE���-0/C�8���<���c����?�yH������W��c���zb�)�: �	ZF���M���l~��r�L����%�Uq��Pgs��R݆5�iJui\��ou��p��`��vU����8S�y������l�;n����I~�%��s��NXrÐ$����zs������bN� ��7\��0��*���荩9w?��:`�����!��ݑ)ழ~�oam��QHެ;� ��ҹQ��I�7�*笽�*��>E��{oc�A�>jO�gY������F�ǈrAh'�{�~�J�h�ӄ�<��M������}��k�Z�U�t���e%k�~ș	��3����W���p��8f��F�	 ��d� ���W�`Uǫ	�a�5i����1-�K�R��5�p%�ӄ��0�M��3W�4��,�:�ɯ
���\q�5;��m�����[�����u>W?��p�|��1ߪu�f��!
b$���	�wuR5nY�g�Ē4W�T����Y��	�%%������_�7cm�:<MY�09�}Y�`I��yr�vګ4���tß�K�v�z�Uj�(�TΊ.�lc�96��>L�����{S@GT�B�0�t�u0Ԝ�- �Ӌ��?`��g��G��q`U?�7�k��2s���K�7H>!E��|P�C�M+��d:���iv1���P(��Q�7Hʗ�f=z�Ѯ�%t����,�;	[����;�'���u�M�pJN�#�&;�A�����r�.�6 �����h�ݵ�~:#"���!�<�U���`�nl�
��z���ۜ��o�OftޕGF����w{J��O)�l�F�kkQ*����oTԼ�b�<�G����H!s�]�F�j�]�4��ΈƸk��|nw��[!���ώA�hH�*�nO���$���@Hq@~����Y�)��=#ZT���P�r��M�2��P�\���L��t�u�L��7
� �r�I`�>���7���W�� ��(x���ˏ���m��r�0�o�"��
|�5��0pY�ZPEŐ>��|l����Z���N	Lg��I���"V�`.���c����"-pK�Q%����b�:i9��)\�D��|�2gu�x��H���5��W�|��;����&���r����?���~��#!�B7�R�͌-W�1�g��D|I���8���`3e�(�+�f�`~=l���Z�8�I�F(�s�[����Dܹ��m�r��h�u�"�kҝTg�8�p��� �R�J-�Fq�#�\��#Ly�����k����S�)��<�d|ئ�)H�[ �������5fjQ �N�Z��d[*<=a��.)�����V��kW;}�XG>G�Ol�Y8�`�������5�T�͹�	}AW��!�y��	���p���<�1��7�M�7�z�1��Ȑ�l�RY����p4I���B�T)�?S��'_�H��"6����o��c����P�N��{��<)�4U<#�rZ/ �H���[��I���?~	�����̓f��Ud,U���D>5qm;� }f�a/G�F�Hi�,��	���gt=��AN�'L/�~Y��1`��P�Zɣ`%��w�����w�^V�T�/�4�Tw[�%��@g2G�9(,K@�,��G4���q���W��z@�\����m��?S�uk��p�B�
���?�5 ��l��� �Ξқk\��vJ�30!��;{�곶�z�L��s\f3g�������;G�֞�&8��CɣG�E�ʪ��kI�� ~<�>,{�8$�O���o6-4�G�>3��ǡJ����hd�7~D��G��w�a�ۅ��R��o��x<$Q�6��Y��&�2�6���ϙI	�a��Q��L�q�^�����q�JX�}��SG�ԛ�x�ּ��Hu�?�/��<$��ĔoK�ݖZ��v���}>�`<�Wc�9��|h��B�f�Ӧ��D��1��b�@(�FbB�bP҆{`Ge<��g�~���S>���� 1XB6F�;+=kT�/X��� �$OlAQK9��.�#,E��Ս'!mj
����{y-y�
���ᘳL�
��q;�F�ך�.C����H������t<Z!h^D垺x�q���	�o9� ����ս3���$��S�d+� Aq��dCA>�Yg�ll`4�h�8��=��FԳ^�SJ�Ͼ����c���Q��q�z��3���X�w�qd3G)����Nt�o������-�?��tC��YB2���5���D�d�۠B��I�S�إ�����2���c^���-���,�������q�nL C]E�I�56�k uL6[�ҽ �#�~���D33 b����t��/HL��g��P�ܛ���V��HP�y@�Fz{-�.��N�y�J#]�(�+� �U`yKP�zܥ�D���}����8�H��)9hH6��;x*{f�p��{Bݼ���|�+N �>�h%R��H������݄Y�%��xX������u#&��R�ʆ���Zr;r�&�h|gY�U�F-q�gl�A���d�m�����oB�@�?���$ojGS�)������y�����A�g��׈��s�;�	��=]M��@���k�Kssn׊�%S�ʫ
�=������ݼ�A4ұZ3�G��#]�ԧ�S���}�E2� 3��$�� H��N�;�a����<��x���w�R)�|��*~������=4�o`�Zֽ�?���N2_�糋�H�@_���u���>��ś��a�E�t��`�#�j�(i� H��L�,��o1*����N����E�/IY���>U1���18Cd��H'.h����P�b?y�I���~ZƢk�r qw����߭r�򄺷�F#�Q�0&~p�Ѹ"kH�۶�޺�jv,ֳE���o�=���4�����%Qq55�Feh��N�I���#�bP6�5c��n�q���kÁ)03yN=�p�3���8j4Z�{����^nwcoK��G$�]�3�J���
�ClW�Q��ph(�(���7<0����-�ᷩ������H�`�3�n0I�����c�3��*�<��%j4xz���R%��e3m$��e���_�|��y��x��`5�������w���m��o�2s���)�^�b{�i �Mo)�j  q6�(꙲�Oq�PՄ7�4��9��K��)��F=�@1�Dܩ�Ȯ�5X��ɵ��3�  %f����4���Z��%��K]���{��ׅ�����Ԏ�yz�>_��"��a�:Ѣҭ �lW����l��nd����7����b��|�R�O5T����+�I� @Tb-�($�,IK�қ���'���_��?�׬� �@����WI.C8ǚ�}��Jl�i���=i���T#�Z����6�~�^ǆ�qFOJ�l� �Y���������w%�4��
����Q~���췇 $^;u��9fC�1���;�_s��~^N4Zw�1Ж��E��<h��W���G����Mae��a�j��#MnPY��/|������l�k��*�j�Ȯ�F!L�#N����'���2�3r�6�����َ��x�9<��Q�``%��f�ׁ�nS��<��P�`�o�M��V-Tu��X�#hVP-���rZT����Kg~�Yc\�~�亅M�P-ޗ�.tcw]�9(1�V�\gHg��d�����1'�\��\Ȧ� ��Wۣ;~���+��Ӌ���E5��r�S�h��Ĝ4e��;,߀r������Z���e�"<Џs�D�G��s��Bz|=�CP)���2A`���xqӓ���y�z4P��z�ihQ&��AB6q��Y衒5$��I@6-7���+AB�V�.�D\z�O��V�G@1����-t���ܡ�����f�pg����?.����\+X����r2�r��������D���A��W*GIU=~���~������Z�H(�����@[(�Yu��,`�;�h�8 `a��*k�9��}�Q���@��#�l(cÉ���%��D��gf�.�'��!RZ��#��y_�ȓ�c𿦒t�|B���t�6rryG�<S ��*I]�ٛf;5(}}�����FU��T��?���h5m1��C��F�N����q���;p_�F(�Ӻ�?����]K7ԇK5;��q@��(ڔ��d-[\i�ō�m���٥�}�K��Z�0%ҋ\E��{�9�.�[��i5�����mQS�3�*)CH�Gd�ip<��ݮ�kJ��e9ާ�Uڗ�~�7��58p�	��.Jt���'������B��J?A�k�Ah?��Q�:t�]��p,goy!�\Ǥ��^�u@�W��3����)��m�"���3�᫩����*6x�@32��/!~w��B�F�:��yyl���͈|�����8$��ᴜ@���)��ɔ���;Q���ć!�i|}����H�U��y�򦀷xE�r����("^��j����\�hE�6����?d��H��5ƕ�[vV8�ʳ�Z�=���m$_�H�m��5 ��t��������9�ȵ�R��Sx
�p��i�b�tr8-��@�F�3�ZBAG�;N����(�����]�e�~N��o��	��k�tb�]ڤ6��<��FP�G[�X����F=��c��o���}V����]�"]z�$�S��gS)(�w}��<� �K�ޗ	�z�ջ'�SG�3;�&pt����E�' �H��ڡP;��g�pu�B�|W�L4
�;�ؗȆoį�,�'q߂f�ѽW$l�$O���;��zǚq����ޜ�!�A��v[33�Hh裵���C_���$%�4��Ҁ�^ɀrfB�{��!�>�1�L&�#(�W�Zy��S�e�kզ��M�Jv|Q �8G~ӥѐI��q��W��9r�����8��` -�c` ������9_�a�X�1H3�F��e���^A?�fE��
�å��r���7ՈzWj �3��93�eé{zh���^o�����Tށ�aIeQS1!-ϷWl�1^Q�:��M&q�;�=/J6�P]2֗���?��"���6���F]˿ᗝl�´Yks�d���S��>��2��L�����K@�<����W��"����V�IQ�Ue8H�8�n�{���+�úQ���xT�����wl�S�e�zuF��^a��5Hl��c��u\��k��{̞����iJN��ce�]��	�ʨ!t�_5�$KH�m;]u[vJ	��?�-n���K���/��@�$�@#'VH��+�5`4��"�fvh�.�O�=��� �m9�^��W"Q�s��m���szbv�����,%���JM�5�5ƻQil0��`rW��}B� V��=���jԂG6%%e�v���T��ϒ�Y�E	I�B՚�����,�`$sE����ł�}S�A��e����`2�I���ݡ/�;��V�c��f4l����ks,P����O$��ĭ}�_��
���9I�����P��z�S�5���rj��j����
����{�PXY7%q��C|(] �a� O�ƀ�8�p�@�'�e�#E�O`�r�[��ވ��˔�C@&g|�i3��#����ʲ ��I�-ښי+0z�6�畚�s�
�R�<�t��>`�Ъ����: �B�10���a]��zfW���,�KP������!o�WH�İ��7��TO�f"�x�7����$fvG4@����Y�GcT�d�4$��9ʩX"��|��	�'������}D�X�8�	/�&�N� �]�?7HD��*�-/�FaaD�"�iK�OU1�`8y�Տ�9�~�	i��=G�k�0v�'�L�qὼ��2ug�-눉*q���N!'�)�EzS:�/��b�`3.��*�r�6�D�ؔR ���GmVi��v_�^S+�6�o�c���� 	`Yw��P�)���\_Ǖ6Vz����;mh�GW�t�]q[����]�C=��)!n\�j��R@�;	��],��/��2gP�K��m��eGn� ���+�+�Ĥ���އV�P�&-<)����a���֧��gߙ�������$��Q{C�X6�6هܓu��1aqZ�����R6��e�I���>6���0을����2�-a���Ȟ W���Z���h"z��f���Jq��I�0�!���\����@o[\:ߍ���av9�i�;m�દW(	\|O�?��t	=S�G������b��0��"��3j��-�xt�e�E�1����m��r���P�B��e�[�f�
-�&\���(�R�ᄒjp�k��nt�~v��F �fjs'��!99�C+�q��?�,5{-'����.	Hc"�<��<��6����`ZK���)�v��O:����{���Zn��̒�c_-$#�Q�A���n�M���hV�7���c+� n�F��gW�/<��E��(��(a=o�P7Ekh�'�7���s��렓�"�G���nƟ��[`y`x^0ʴ�1��݌���~"�M�l��׶�C�[����{9�p�����]�~�:-98���
�}5����~3Z�G�]`}��?���]��,	�����������VAym��z���=��˦.E�Y~�π;�G��x'|��ʨhҕ~���){��e(���rLW�|̯�ͽ�N�h-�0�09Rd�;u�+�O7�	�UT����/� ��Cz��@4O߲���]*�;�K�vO=_&@�H�3�����dtIO�'�F-)�$V�v�v�x(���u�o�ue]�sa�{�M,����gd��U`G�!��b�抖�܌��w�ͮ�*��6&��g��_��H�`kR�`�f���!�dيK�R��ᄪR��K�6o8d���%|�G���Q��oK:����t;��N�+I	��[i��o���(
w���ߦ��Hf�.֝��r��1{�=3��
���R�6�� �l�!;�W�Ґ]�t1�O7��������#�S'���*F
��$���`�ɓ-�Q�8}�jo���d����E��_�m��n롻�Hz_"A���D0�g�[�%#
7%�洷�������|9���8�3X�%n��ֺUIVo��Eu!��p
0R̀�b�)tRtf�����_�v��^w�k�o���Z:ʇ)����J2�Fגta(����)�;4k{�:�^[ny^u�-B[�R�
�T��b�F�r?�z6�F�ajm�5KH�����1�+m7��xf~�A���'�]�g�[�����VO*O[Ε'�U��J�O?	�u/a7lO�}�6>p��6Kg����9�?g�i?�2�&>�.��4NJ��!��G���R�;�
�%� '$�����m ����k1ݧ�����8��O�K19�8���k���7
 ��!2�V�y�{�u91_���*�*ϖ}"������4iM��t>P�Cw���R��!�8������B(D^\���Q[��T�h\�s֔�er$jEߧ ��Տd��6�|�5��f��7t��"E�J ���5f���V��,�ず|��S�t׹���i"/��l�p4��^W�a|)!ʸ�85�p���͓m+�U^��qc����dy�w���(1g���RF�J�A�(�v�X���:��]��X�Nm+о��&Z�l+AY6*���޼zl�iw�Bd���Y(�3E�B
,��@�	�p�z�|�d�L$fs �ߣ�*ZXNg��ڽ�!�z=���ܜ�f��htp�ْT�Q��Y!�	o��r�?#�0^��Ede�­�̀��ɫ�������'sjQ�p�w����l7{��B��Jvf�do2��$qJ�ɇR@ҶO�MK�OA��&`�O;�È��@"k����4�5$ �g�T�x�G��V�ņ2��z����V9�����'���5r���nc+�q#y��>L��'`i�j�
�j�¦���&jU�.��&��)F�u�����Z��L�%�m�u �{�xE_S�0?b��k�d1���0���d�xm�a��_Q��n�|�B�;Xcf�]�7�FjO�gٻ�e-�L��@%𪅤^ �a�@[U����ə����R�)��s�9\fQ�̾�����͛v�BoZ��I7:�=pSи����'��]p���hʁ��q8r1p��"��k��O���i[�n�s�nb���j��_6�����7c˧$�~ԡҦk��8��F�m����,k����ް=����^揫N�r�O[��i��*nL.��o{��s���?X��sz��?�u��ݓ����>�Z|��D��z��
zd�m�2���z���>��z�nM0rC��7�#|4'��o���L��}�w�ʤ%Έ��D#�ac]����.�U=�J6��R��T�20�"�� 7'�đ�
q����iQ�RzZ��`4��3'���XfS����c�>X�����i��F>#2A)+S�g����H�b �U��+Wc�0v��a{g�yJ.��c/��<�G,+D3������S�Rq�ϣ���ږ��A�}�g�3^2ٖ�0�j�=2RG��f������l�̙*JHQ����8 �_݌v��:怰!ʓ�Y�;ȭ�|UI�&�4�k��1c��r��r�?4��E�P;5h���.��(��B@�H����x�oK�b���S'�k���A&�Gx�*(�8�NQ��NpI�|A>GH28L����mN��Z�����j@�q��:/S�n	�cqQ��/Ϸb��i���j=���ƒ��$���0hq��	F�w_wr<�U/�r�J`p�WE���8`<	2ӕ�/�v�'���tVU�&�C����>)�j<�����+b�;���B�1�pZ��J��������٫�.E�]�����q����������\4�/l3�t	()Y��+�y>ʯnb�Ļ^�P�{�"�� ���7��:d�
� �5��u��8S�x��V���M�N���Ib0�KBr�E�>� e\Q��ټ�2f��@�cFI�Yz�'ԁ��+��{�yVk�4��8Y:6��1|��0��s�T�"T1�ƫ��<�CȐ�3�A�p�ɚz��^���ռ�bTDe�����.�1�V��D��^��`H�V:VH�4�{���/�K��1\� :�7���檴��]U���+�w��~;ܽ�9�HC�|���.K������.��'��ɔ�Z�7a�/���<�}�)�&B��>��7���~�f�E~���6�Hs ��ڶ��.yF��U�ˬ��7x}����ѡ��v�%`r�LnI(1����hd�1�_���ݡdu��%��	d��&O�e�/��Iݱ�l�r�R�hE�tW�Y����\K���Gn��d����Ș�n�Q:la�:�{��r����
��%��	�"{��n*�I�ڵd���(��q܏+ZZ`�s3|�m��8��tߊG`p)�X�bJ�e�#|U��K��Zn��`�Sx�_\��V�=p��3y1h���;F�`p��^D _���LOM:p�)M!�~#�c5J!PFOJ� �O��(��:1���� m�Wi�<!�̈́h�D«�ϴ ,Z�ZЮÑ��CQތ�s3�P|����i*�#�
_���<-
�e�hl6![Z��)��~�����Q�,�!.t�Sͻ�n�%��q�ʉX*{���^���(Π����1��JP!�q�x�Pڊ��*���DB�6S;b��)D���'��̞���Y�[
Ok��C�H�a!�D u9 œ�3���, ;�`H��'�aj��Ш-Ջ	k�N�,��U����Q����������V�|�]�[�����1�٤�d��sSe�+��ESz^N�E�R/7�q��ňk�crGR	������g�<|ZF�ș�
�U"\D�sD�l��/N���<�M���IO�a�������.��$���Z�k����V�T�>*�ٛ�����C���`�EV��?�k����E����������~J�a8�(��[������~�o�Ɗ��R�kj�Y�Cr_B�f�]���U9�҅���{2ݲ�{�bn�]s�E�8u�O�Cx��V(�FV�e]� ���:�Ɔ�6G�
�py�E�&B�뷮��{��f�Z㚥۬���X�5?@�}3��\ob3I��k�d���2�\��x�F�v��эoժ�3�u�3Io���~�pM�;�"K�W����s�Xz�R8Š��a����5���|.��B���j��"��9��Hqzx��v�/�o9vd��Y��.o�:�����:�=�Q0T����St_�#�w4B4�&��z�@�* �C�|p$U���Y��-t'��o��?�/R� u�R./p����:��������t��{��:[�HU��ػ:bcC��b=����J�g$$@�)�X��\?�����P�a�|��v��<2*_G"�I������I'�`�j��������[A*� ��M2B$��(Dx*w�~K������q�m���>�
N�u������wv,�	.+�Fxޤ��fjk���~w�<&ɤ�]Z�t�����]~/��щG�
{Xv�Q�[_���O�Cf��3�܍4�I�xZ�"aR":^�8�����z���%R�(C�v5�"�Ot#3:��{Zy$fݠ��Y��Y�~��B\�s>�q�Ng�_���Q��ڕ=
�R{�0$�>���m�^AaDg�q}-��{�@r�o)n'I��d2����}��c��@BZ����{���z$(����!Y�-ӛ�&xٳ79�nb*�ǈ��F�I�pC�0����F�qܰ��-�
8�	�W �k�&o��"��#�qs�TH��sCO�'~��m����G��=�	�����d�:�Ѐn���fx�>�~P�m��W��t's�5aU��:YV;�g�S%l��h�pu��+���W�E3̧����\�]<O1��fm�{�����vkLl���L�W�U�����w|.;�v.f�y�B�/�a���y���V:��z���X��'ſZ7o�N	_y7��j<m� ��P�ѣ^o.7�0Q�EJ�hرS���W�}���b�	�$�E��-�9�_�-�eu���tqvRN=�;1��KF�#��I2B'���P���jI��@�I�B�)�]c5Z��;g=��)����p�R�ZTf�J�\�u邊����BW�hĶ�~�$ ����#���AV��g���X,��sJ͛@��HEǛ/��se��넙}�%�~��v���X�� (��ɉXS@ٱx�?�����S{���2�RU#� �����)ZQi���_�U�B�=���!�Ma^�<ǲ�(>�e�(���	!���P�8�P}�'��^g�$�D$�:̾�\���Cu�TM��~*`�s�|Q�ź(�V�|v��M`D{���;r�����-&e�.<Wq��GVK����2�#��.�@�U�gf��[O���L�M�=��f��aM&x��R\�!���ޙ��C�#�	�/[PM��rq�Zx��[s�r�CX8�w�Ub�R�{��WX-0H:���6,������[�PέB*���<9| N8\��~Ns�t��g���Tt���:����6e�l���&����w��{�4�V�z��9.�-P�`��g����i����=��&Ŧ�0X].�$KvS�6�AH�t?�s���	������]$-9�HP��j���x�!�nX�{�=E�쏩Q�#$�!1��a���}i�nx� ���M��X�9*�
��#�  �W�ta�Ư��U� [���
	�wp���߅mCr]I
��jS�;K�*�X������<.5����q"��VZ� ��0E�A�{�;S��jV��BlٱK�?� F���'\[��=o���7�j|3���\��4-�EH:���	�7���b��w��]����6�1�4�-����5�-#wq!%`�:����8M������a"�&�λ�VD��)T�o�;_�B�t �X��NA�꣦���W����~pgy�8Ϝ��{�ԁ'���f���]�A�_ίjJ�(
2iL���py�����0a���x������G����sO�F�xl�I�$�ÉtG>�,�k���~�?�F����Q�^�:G�5�)ʧŁ^�9���:�1F��Kg5����q��� 5gn�y*�d[`pM}�����ʁ�T��F��.���qR�!n�?��t�U��Ŀ�3� �B���ji��?�����ؗuj�٢?���0X��yj�[�_�W��R�� �#�@��D�7���Zn5�*Cm� ��d��*mѱ��4 }o�hm�0p@#_"�9I�n̔a����ķ3v�k�`cPW�U���!�U�$b��A<�±Ŭ�+�7�_�MqYc,�v�t6�B�~�tQH�'���`��K�VN֟�#C2!����!_�-"�0ď���Wy*Aڵ���AOK�Lş�״�2���k/`���JF�L˴GSAm�tFA�2��-pp�B��(��A9���]��Y,�ٓXWQ5�$�����P����4�X��,����B6�]�Z��Io�&��u;�^�,H��Gv�A���
��=����
���Z�*���$��A�&���g�mk�4�m��)Fѽ�K�{�>Nɯ,�G�g���?�t�����؏`��)�A�c��=���"J�d�©��p�vq�_s�%��y�W��ʽ���l"�>p��&|�.�fg%Ԭ���Y�=�?/��~ m�_��[w�:TI���/��LY�7�����_�����+��e����R�vH�f����*\���j�x����i�g���_�����z�$�̊:y��XWW�|GZok�kiɼ_ݲO�jR�R7����%�st���*��;D@dT�:����;I^���2����;^�r?���dD9����q��ST�ު�S����]��s_nb0¨�'��.�v�\"��1�j�fw}QbE4$��q����H��?�j��Jj���.�Dru�N+�^FU�S��D	�=�{�4J�,8	����p�Q�o ��Qv���Grb�bWMi��'�����t�<8j�e����,F�,�F�Bn�,�.!�����^����Ģ����S��H�ѐ�&��8�Q�V^R���Eǡ�݌ˠ�Zя*N�5'Z�?N70�r�S%��ьQ���i�ͪ��E�*{�r(h��D.�t�xc��kB5�O4gt�"�����(!���BTkA�X����K�V�"{�*:^�N����"_��,U\�J���Eűbt�'g�L��w��h&��x�LB5maBG�����])�:u� :������3�4bى�,����8�
�B��n� ����������-�6�jem?���$ղg�*`�Y��^������1��̎�zr���}�,D��).[I�^A����T������+Ta�%��[l��m1�i՛��C+f>S7�=e������G���Y�.�����R�5c<iw{�Wc��W4dklwqg��vR=U��t��a3�}�O�/��AG��5%��hW�#����T�	��a}�pɭr����e������#C_o���b�`�Uy��R�������cI�����C�4gž��i�.{�3{��YN�!M7aG'Dz���O��I��c�.�\G�R������w��`m�>;7 P�{~��rH�7*ԍ<���童�,=�u:S���>?>⚋S�������Bl)��0\H9{93)ϩ���	�X��h%G1���t�=���{Te�a�ռ�*c���k�{lNy%'e��� ��e$8b�.��1~۱���c�q$p"r\eso�E-��������..���ZXŋ�<^5�8EC!=:��[���,M�jή|�K5|@Zv<�_ȥ��c(��|2�*)�6IM�v|$3k��PH�� �0�3%��^��ƀ_��ܛ�ؾK�s:�q���(}�L��>�W	Q�#[�g\%���;]�x�8�ԯ�ٷ��?�:#���m�e����&������ɡ1A�ڍ��$��˘*�^�+r���qH�Z� 6���z�|9\�)7r���K����ս�{n�&B��uܩ�s�F��T&M�/�C��Lq�ͻx���u��|�M#��}�̧yV��$*5��pʓe�.fu}GS��)IGG��A�p27��]�ΰa�r�D�'\!��o�k&5$�rK3>��t��"l�c�L�Ջ�\?��7�]�6���0�p�ME�)ޏ�ô��L|m�ݒ���M ~����r*��7�k��]�->8k�A�td��j>i��ux���"0�# ����(E���%h��އ��N]�x�F���	�ʜ��s[����ħj�LU�9W��D�lR��Zg�"���)7��S��0����[�Vh t�氓��{���a�>��2%����;�Q����1Ba�������lSc�z�[r	������<~֥�1����&cp!V�p�����^e|g#8��?��Bm@ ��:n�$���3r`��}vD�IuCi�A>��*�@F@����뿙�o���߇�̵�'�f��HۊQ��.&��n?���Km�<��z6C�.�K�e��ᳲ�)of�p� �(�(��YC1dL0ei�v����(y
��k�ǖ�Ӂ�{��iy��O�R�ċ�52��A�yB`���KUC��PR��U���&�m/�2,�s3*�*�_ ���x�e�i��-�("n���w�;�L�/���M�JFKP�"ZU9�)�>ֶφ�� ,��"(gܵ�J=�������*.�Ev��!
�����
}�o��dYۆ���pCI+��V٫Y�M�+`��?W�ddn6'7��|����L��.��Z����3�YoƱ�J㠋�(������qw�J�-x���26p�P�Hp+�B3��L����DV�BO��ȏ��.�[$��Yy����q�ʭ�q;����`��!�N0�x�
���;`K�/����5[
;fL��V���l$�ٲ�n;�کiʌ�j�ō���;z9��h1!?@��OY��@:Sb���o�<����z��$��'clcG�$.�En�Pm����?�h<�@t;�W��A ���\�ô�����}�&�Vjk�Sw��o��(�/�%����E��I���K�S5�Z��dJG!�V���SRɄ�D\A6:��
��X������8����p��♚5FK�� S\�F�V�c�X�/ũ�S[�
���~�/��v��#���{,}8J>t��]��U����m����hb�K�Y�4%KƞO�4h�2��d��ڕ ����dtE.*9cJ���q�X�TQ07�D�ӕ��)ں�u����e� �+{BUJ�v�H����?g"Ʒ��@���|�����n�洈�:F�e��x�ܠV�j��jn{�����Y����ȧP�������RX�L�F�����s�aAe{�	C�W�|N�fh^�������.��a�u`�:����e"��q"ab:���1��T�8F5u��2p��l.�Lz�EFl�#q;�
�g�$eĘ�.�h�EU�s�ôv�f���9K��z�����f�J;ݳo?�s��nD����R�r���?���AxQF) w,��dha�爣o�C&FI��&(�0h�>�Zx(ۤb����ڧ0����RU����y<�g\����|���R7u�s��!ߏ��]Z��n�o��4㹚3[���h���.Ds,h��K�_�2_�@Q8T��2� @α�i�~���-H��zBI���w����`���'d�O����T>~0L��!�򼐑�I�!�Kr�HN\6��b<�a��ewy%�e��p���Z���L	.P�K&�R��SYM�:���
����Q)�M0oQ�}�Vt��Q�K'ј��b�9�;�u�\��%[�i�-g�d*RV˶���x��c[��Ъ��}XZL��E�?i���p8�/�
6�bǴ�������>.~,��o�0}�B���Ѝ�� e^�vѺ��r�p��9B i�}�-G'W��8�6ҩUW�j�����5ʊ�`M�q�@FԏS{��$v�N�Vo\ӢqZw��*����g��r�Cr�k�_��jy�	,:�0%���ehn%��WT�>��Z��6)����k5�������ᆩ��V��a��5�7#?M�ZτN����Ŵ�E��nU��H���+��Dhë�o�P�φJ>�,"�(#�a'ѰJq8΍��Ԅ�N��<`�ށd��e�&3��d�(l��뺜⟨��0Ǣvzկ�� �YI_��V(�k�y��q�gzf�z�����[$�A<ڴ���&R���;^�?�+��Z>΃�P��qI[��q�l�\�ǿ-�S�AY7�,�P����rC�W>"gW%:^��Iq>S_h���5Y[�Klc�Wf�%kr��An�l�^J��r.Ol#��^����ٖ%웄C�^߈C�/Y����> �;snH���	�"[��9  �?p�l�p�B�_�͘lNb'H�:��1� ����dmȴߥ�D_���F�Qj��Ċi�y��^ �+�ڿo���J�a}`�[Z5�H~��З�MW���'[�(W�~9�A��歑�����}Dq�Èx���O0Z�)�;1'��q�v۫۲U<P���#'�']o9!w�}�}DH�y�e���(�;׾��l�:`YYd��&71�]R�����M�$��FW�M�p��Tq�eΗ�~�H�lń�:�!١���t�^��^��۪�`L��'����ql�v�É}���������y���ϝ@;�0N��L$!��"�u[
ZgU��Z��_�QC�����{J7�
�lx�E1�Và�� $�kmW��_���6^i�o�KXT$�Qz�1�)���6tq���o)h�r)&%ڏm+�g� nd�����G4�z�Y��8�aF,�5�&J�
�|�M`��`җ��i�0'"�r�*Wŷ`OKx�u5�T��;�p��ZƔZa���i��X�'�X�!M� xr��M�A���W��ouOk������<��a�f����w7x�d~ˊTf�G�h}���`Hn�[;����g��
�?���?���Os��nB�qg�6��������pIaP+��ȋ����3>���/ېT%��SZo�_\8�y����Ī3�����+Km�\T�=#���M�,0�y���ʯ�M5��p̐H/�9ga������9I5�1���R*hH1�0la��J���:1C8mw�g�����\!��彝�
^����i��<0hL}7rY�Q@+�=���2�
=�g;��bT���"PC��������g!\iv�3>b~C�`^�,V��N6=n��U �p��x+g7���FS����ai��&b�4���!��i�C���Z4ʗ+Cp����ķIX�� $(�p�,U��r�^AK|���̋��)�1���D1g=�����!sl������	9M����8��fػ��k�q}E�y',b�0s�G3�4TR"��~0iF՝�����]Skp�p�����A��a��9
1-���F;�!��U�c��b�] F�b�e�ڔo��J��x:=u)��+p5�=��'{4��w�p}KsS�O�|���P���9���_"5���:��mc�e�t�q+��>WzO2/$�R��$4����XȤO�`�烡������E+��i�]ؾmVZO,P,"����z�Ʒ8���o��v�Z�}?�.Ѳॊ$vl�{��\r�,����'�J7�ʈ��m����)�i�4��n��5�Հ�������Iq�8ճ���V�����o['K
��ty�X\��F�}\�E���rW�}va<5���$�/9b�R���	+�@�8���u�N���7���?�C�^[�Ro���\y7�gB���}*f���g�hf_P��*5˞����V��2���L�2A ��9�'b���:�w�]�	dڵb>r�Պ�h|ea7��jo�T���Q�-�G�����C1�L(�(c_�Q�8f*r�N9P���{�d����a�b�5��d�̳\�N6�#S���_s�2Z6�6�჋2I@#�j���my�k(ppw�̈a��,|:�כ?@��G������I!kS��׮��:b��"(r��x|�_��w=�&�\�Ӻ�R�Բl���We�Gt�`({Ѽ��M8�G2����A5�W������ˬ�k���q�Uhq��P|�(�'KW�^$z�=�%�}�R��7t'�Q�`ԧ��B>���e�F��`ivX^��o��P"dľ��^���:��7��[�,��
�ǣ$����rQ�G�,�xQD�A����Qŏ�������q�A0ETt�a[�2��<�0�a�,S�ei�i���+��@kTQx��Dr%�����.�\匿�l��Ƿ��/K��lpL�l<t��J�����q�S1�>S�O$,^Q�����YE�Dˁk|K�QE��@�K��o\�ȍ��t��8B�'��8�t�V)�I�&Y�	MF�7ū�ˡv[�i���4; |�Z.��������X���ᬨ��� b�������v�v��K�;W���t�=6�%0��+��K�j49�����t�2�ߥ��&E���j(J�t�Q��?���\�fG�Վ�
~'$3VY�L�}��F$�q���jxX�r�����}��!8��1�1U<8��^V��kSo�/�䜽�r1s��`������ҕW1#A�K��]���S.���G2R�s�N��</��ŬH���1�Ƴ׎ew�+"�>+ё��/Vt�f�x+pf*���	0�{jD��2��K� ����&��$D�m�	KaJ���$K�'s?�Q��N'���-{i����)�HhO���* �����/�C/p��=�X4F<P< ��� ABoP��q)�r(��$Q�>�������4�+?�LQ�=����ש� �Rwk��^dU���#J|\��R�Ug�q��%>S7O��	���Jy��8�f��|l�?�����!�cˈ!��X�F%���{S��N�^�'�ܐ\��}��5��#��]լ�t�W��:yX�}q@�]��8pOu��j���$����(,j���r����E"��>T�l%�Z[X=�|�%�2��J�1���ѓ�4\�$T-2�g����,:F
:/�ֻ�U�2})֊���Uf$�Ȣp)��}�m�����T��u�h��m�>�����R.+�Ee��w}�����%�#Y�	/j$�C�߼��S��*�:�� d,��_�s��Gv�?��dSp��܆آ%��-����ٳ06S�+p������r|�� -��H^^Rh��d�<�=�Nvg9��_��ᥥ�h�u�eJ�|a��$#6RU8|���!��>��B��Ax���
C&\쉯zSυ���j@j�ᒎd���B%�����d�!�e��������B�+�E����9D��<��m�����z,�{S�[�ó��}�YI"���,����`�� ��NkZ�в���	����Q��-�G\��	_�8b62r�5ܿa����������@kh�����x�7��27���C�V��c�����>J�Gzg��R�R�zO�6�!T$1�]m6rL��*���a��W\�w���i�I46�����CB��F�-E�/���i��2.�=D��N�d�W��JҨ	a��]�`�BpbSJ���Q����������f5�]�L��t֙���e��0(����[�8�Y~�4k���\�j�˚O`'�,����������I���?A����N���)�q�Ņ_�c֎D֓�3�ѡ��� ��Q�E�g��\����r���BmȊx�܊�� ���õe�"�,�͏��k
9l._ ��P}Dw�k�	�&A���+CW�Udt�\�Шb��_��DxU9�������3HE�w��G�����Ԙu	��!��e/���8���oz��hd~\��
�䱣����{/[4���+�@��ԋ�^����,�j�6�}eΒ�[
�R��r�TE�������U1�=c5��!5�#5�fO�`;�n�,WP?����������9�����9���086��
p75���r��=�^�D��ki�I�|�^�1ѥ̎Op˾���+�7�l1"[G��#S�'d�ɉE�;��V����-���ōV�#��c��(�ɥym4��$`�.���2�uw+2f��r��J��T�^����q�⇜O���?�L\*.�6��@�:�59����$����Z��N-�)�w���W�aAͅ:e�0�ם�5���w�e��b���mγAp��VY��l ����/M��P��1R�g㬦�|y;ۑ>n�@P�_Ҽ���uOn�dWދ1�ZJU@��:\d�`Lx5<�����<��;���N�Uk�
UY�qE���,��$���(?�Y�?p�6^���eS��V�PW:�-�|S�)ڽ�JNZ���lT�q���e�B�`�S�o��Š72���ы�ph��|˖=���]�I�d������_P�Q[�䀷
]�����9*�9I����u�� �'B����6��x�si�z��s�4_���C������[_g��c�NUBIU�8�b�őbTF\���~�!�[g�'[<��5A&�X��!����%��B��M�����1%;j����Q��+<�HXm֊�=�au���3�A���6�����U)�0��Bn���xG�\M�H[
%4�gi�� [�Rޖ��)Hi�P��+2��p|��@��ϴ���e���	��Y��i�8�0]�k!����O��rUW3?/P��"��\��G�oY�ٻ��i����'�nDѽ�VEH�!�
s�	�]�Ǩ����ʝ����ީ�e�ϜR�K�*+� �*�W_��nR����Z�����D�J��7k��}?^�Y�E���a��{_#��� �ZY^�� nR�e������ [x�w�Xy�����G@KU�_�A��W0��\��P��T�_Ϡ������������ �H��p`:xGR,!'��c�Ƌ5�4����0�$<�W�D6���(JD��l���)Z*n%2��#�������=�n�r��*������}K�q͜0����hBr��#���L�P������;��g��E`$��ve_��*��e�]��W;o��*�wO<HB5I����2��;�1�+)��iS��L�	rż1$W<�ƙ݁P���X�#��&�횵��F����84B��{+�p���a/�1F��qE
&z�a�J���Q4?ȣ��"���>�#�77�]b~|T�����,���s�>-ո�ဳ�� �<8���8J��.��/`��ٱ��}�S�aT���x�e�{>��n�� ��0F���Y�ؓ�i`~S\�S��&��T!Mk��2UY�	w<!� �� 3�b�)�	ͳ|"ί���U�pj`oB���@t��R�x�|ڠ҉���VЎB� �(�X�uT�K�`/�Y�~K��a�*ڣ�s��:8����}� ����K`lz�x�XAQ6�lԣV.�-�a�10L kt� ��y���z�/\�M.^�w��A$�DSK���"�%S���� 1{��@J�}�.`�*`OI�W�v�q��I�@s9|z�0��v�D�@�~g��E#�wM���iAp���u�`$�5�٥�[!�5�F��#�� �z9���!-	����O꧆D���O,�"�1s~��H�BI����/� �H��e�JvO��Z�{,ET����a�N�4�>N�0(�[%�~-�:ZɃ�$N+����`�);3�K��Ω\������J�:y��ԓ��j�q[�×���m�]�*�c��u���>s�/�{�P��*�B�T-�������{�۔�N�w�be-�LF�Bң��4��ET�D�'��?�l�.[��66��6@��@M�̓a �V`�5n��%^�G�4��,�d�
���P�u�Z�=�G���[�6(����ta����H���<����A�����ޮ_�QE�|ք+�T�S��4�΂�%�&r����������e������EF�-�b�G�c%�Į�#����}R�"fH�2ې.�}�~Ļ�z����	��S�G��36d�s�BDc\Q`�_���A�F�n��宀�
�)�^,1J�M/�X'���2&Ѳ����?��+�#,b�P` ��"��J��)�B���8���7�wz?(7�	ҹ�HqR��ւRsW�x�!ʂM*�r�_~�WqS�v�շ�$(%��Y�sx�ҿd��A�]�wYr־F�0 #*�G�C��=��)n�(�E�����,ԁVȞ���&Z����mՋ���m$��-���F�ŁZb\��D��z�G�n�QY�a�V�����/y���yX��H������m��M@�Q��jFXF�tFxҨДxZ���| �� ��C@OUks!j���ϵa��h��#4?���D�z�mFb��}�'86��[��<����j��V��F��h�z��-պ=�~����U��������ŃAZ����rb�gv�nu�]>bkg�IARǕz�٧}+�!�y�ţ%����C���<�T�`�~�jF�9��LS�����BC��JA}}"r���- ���4����W Bn��m�����)��mKN�F �Lh�9�6���� �=.���4���a�X�=c�f4pƀS����x�Њ���Ǉ�>J�תMl��f/;��C�]a�8��h.�dN��M�����_\4,�R�Zn0�'�TΏ|�����mM��tH+����g�������ر3�G��g���Ti�ݿ�
YH� b����SuK�?�c�Y�P{�z;
#��>j��Ȯ�Tw��J���h��5�]f)9YP܄L�zX-�uq���d2�ʟ&�آ�'�ԫ/�i�AD��2r �LQ�Z���ڞ�pM��˷.�m�u�2���°w����xQ|���/s}9�x�'YoEuf�/C����$}�{�d}�Ya���e��r�I�M�|GqH��2s$��rFhQ����Ky��^�b%��VW�ߤ.��=׈s��b��<#�� V��֡���ڵ�c����F���*;K����*�7���츤���޽XT�<�Ȉ�E!��Y��Q��7�B����1M�\�m��Z���f����7	)=�m��ݚ�~��b�p���\[߇t~�k=���S��e�/a�}�"�d'`Jx��J>�/�P�W+�Vwd��N�~w,��1�I�~���"���r��ς��,+[+�eѰe�J�̰����@ysA|���y����VW�8�7�ى{����P����@��1�f1	(�"�LvT�����\��e6���-D���-�Gztٸԁ����˯	2}�'֧[ʘP���Q���M�U����_������9Ģ�ǫEd�u�֚�:k��em�"���-�����ܶ=X� ��¶�B������Y�u�[
Ho�Ǫ3�M4N4錅��c/<l?��1$ϯ��S��:8�/Ri 1Խo������mW��߰����.�����X�WW@���_�[���~��͇�#�S�"�/��["�A��e�bW��?�;�s� �Q�Z$�*L�?�����]��"��
yΏ��e
P�/��1J�Ů��5D�	}�U��,�{{;Lz�|	_��N��7��� o�6����ˢ~1��`nM����O\�A2S处�҃;�dI��qm������� �d@��+�^A� ��	��~��|�A�ZU��2XSx~A)ef�� *1��H�����ȕ�n���V���o�����+S��a��D���bھ�E#/�l^ W�s%8*���ԉ�]�t��m�Fy~��V5n��Wݤh�"GZC.$/��W�xg9��.��O�Y��76PG�E�I&��ȉh��-ߴ�I�qq/!=U9ѧ����thm�^@d�&��:��a<����Lߌ{���pI$|"�SsC�]�-H���J����S�\��/��� ?@E'C�Go"d{۰��ݴ_C�՞#�^1��ƜN��1��8d�]��Y�8Z$��?�/S�1�xH}6W^
LH�p��C8>J���:��][��s�`��'�U�����!�[��Վ���R+�vqn��724>���l��x�.M�HukTݛ��l���m���K�C��b���-q̟���l��6�y���t(jw����'���ڼH�Xj�w�6���NZ_F�����7-�&����IFZ�<;�~�xM�u�H8�i�7W.�|F"(���f�������S]��I��<tÎ��%�E�V�N��|�:�d����	��a�Di%Ѩ$���9:̙��ᚶ�J���w��r�zG�7�%�V����'��ݮ����׉@�Z��R�������G��6�B���jQ���KE).W-�{��Ӕ���J���h/�6���
.�	�Q�,4	��bޏy�*k9A���p�n"~����sb��b�;-4\-g������Eݯ�j�>�߮i�ݔY k�sv�hޔ �s�D�5V�i^+��.�Rf,�\�D5�/?�y(�<�ݩ�:Q�@��[�׫Wr8��C�H)���p�'�>b�2ebv�j�v�3��x�5�5_R���B�6v�Ԗ��*d��k@�X��]M$�(�q`� �����O���lC-�rK���j���c�����uTQ!��&��D����ȳ��]F�۹��3�'[�Z�K�Fi��\������w���q��	�9�c�g�a��6��*>men}��j��ˈ PoR~Lsn��
��.b ����S4�?�2��_��+X-� q�C:�m�
��adI�f�1�|+�"H-�ocR������ZX�X��wi���B Pu�!V[����0�@@�����$N�wt`���f�\sdH�i�j��Ҡ�&�l�ǔi�?��ʶB�TKPOҋms_��,�=+�����
�z��7�|���,�=�Kߝ���s�#l���:{�!tX��[?�$N-��I�Q�j"�ͥ_=��sR/�;���T�r4G�6"m����gb&�?7&>ݣ{D�gC�� 1�icG	v�OC�)k��t'r5���L*%�=L�1�|Լ5��л����V���K1���	pk�!Z��3���E���]!w�G���p�@3��ЙѸ	�K��B�>����X%�n�3�����B��o���3��A	� _uW!�=S �(
�8Q��	
�Q�^���;:�O�œU�i��r����I��c�sR��>��;.dp���x�iW4�i_�$|�!>�l���Pwc�DG�C��	"(�r_LFH�Ga�.`�u88NP�[�U>s��T��^Bs�h���O�� ���!ny�2۠�Q����W�O�UM����t�yV4�'ۺL2�P4(�'J2�":�r�	�����ĹK#hN˗�I0�z�s}[N��dD�t�$��3ɲ�pD�3z�AW��_�/㽞ۤ�>�O��#�E��9�(��9�I�7q��8O����x��+-n�L�Hݖ�'�0k��D�x/^OuN[�%v��`����Mz�ø�R�V1 ��wo)�[�|k
���uQ\����{�A�X�E��(܎H���2�&��h��"����{�t�p������$0X|�+#vC�0e���Mx>��:ۈy֧I8 �SJĥܸʣet�y���ɾ���-ڊG/�nx2]M7�p2p�?��{����(���wxb4(��:�6�0����nv�. ��oS�ǅmK�q�]��<����������1 �=�����A�� ��S�5�K�L4�o�M���0n�� ���yEȜs��Cm��Y�K�Q�rx��E]��J���@�]�����k-�FM��v����(�=��a>/ݕ]0�21��=��h�=*xs�;_�h�X{h4���P�������ta��&����Y�BvH:ފDS3Ă<ҍh��{�8��g����%+Ƽ�p���C�%"�WjcM�#!�z`Y�E�J�V�_��Ì(ua�����F�ƛQ:�U@��%je�U�q��� �sձ�S���[<&�5 ��(n'��k7Ci���J <���q~WB�jl�_���r�,�۴϶i��l�)#�-U�W(G��Ц5�T�T}�@��h!?T3J0�1���`r=�-�bBT�Θ�o��t�z���>Q������I릳�P����C3l���(�ѓ\���0Ɋ��̽-ϼ�7�z�oPk~��_�Ѹ�E�qfS\6��U9g� �*g؍�+���E���8��zAQ�� P6�qc���z:��� 8QD�$�㤛��w�� 8���fnyz��0�j�_cۄO[���.gnO�lEZ9{�&�1�ʫu8�Kz�l��L/w{~t����JZ�6~��"��cg�|���L��� ��+BKH�EF��U"�gV�&�����G��/G�����"1�*��!���M��T�z�:;Xf�x�2���T`��S{�M��ʒ1���?>��{���#��	�]I��l��Z���_a�[��(��e�qO�	-m�7BM3���=�/Vf�-�/��7�J�e�4+�� m�=�{�y`s@��$AFb�_���M]%����+e�R|�_v����O�ibp�1|�+G�sH�g�2G��B4�F#���-'�e:��r��i��a�FIẄ�Ͽ�c=�מ�NzI�h�+]��j")�u��x����U;3*ҹ����T3��؊��v��Us敟�r���d��spp-��(n^���6��E��|.��:}ՆL,S�n6r=K+y���m���	d�����]`r�Q�\��7��/��=pŵ�Ά� �_�c��dPS�E�1������n�e�Z/�I�a�U��
�w�5��'��o
VB�N���*��Z�ǧ������	�.�SYX��ǒ\T�����ۡ�5ظ�k��]���O�+D���bN��~v����[Sx)�+��]k@IQ���H����'�&9pQS���h��f9�)��<.*H�M,��Q��.��f_	I��e�RJN|B�~!�Q��������U��Vw�^�Q������]O�1��q\Am�]=ѠMq*!�w��O��~0"�۪�ʨ�q��K]lV��'[:���P�N�ֹ�ӑcTrq�$�ޅ�G�.�[D����I���cض�lo�2�Cwr��ϙ��*��G� Ee���� �Z�������j�56;x�nە�8Oj���y���|zvo�p���i] ��jw��sk_n�b��Fʉ�#�G+�?k�a�H�sb:��ȃ�R��ơ����� >e�ip�Lk0��ȘSޤm��Z;��b��b^
�i�����vrV�R[Oi���]y��1������j�C���&��Ȯ̝=Ij3�T�k��*(�-���' � :ACb��3	�EB�dr�L�"���SAA �0`HLU�aoCE6��s���h��6��}���֢�D���T%�	1���=���'R�m��fcT��|\\�L�X`�lV�-M݃.��A��3X%n�g&�������Ztg06y����c���=�1l�~�01E`�-�f� ��|�Q�D񊽍})��\fh&�t;�<Л���Z�#ij�����4T�H���!J�M���2v��4D�)g��_���9f��b-{���R<��Js�d�p`VG���
��WFۗ���T�rА��Ex睽��Jn񩋪C����h���>��x��T��(S�/2@_�+�X�f/
�&"��n3ʲD�� y�Ѭa;�QG�Ua���N�#�8���ڂ���ώ�Z�����u��U�DB3��_8��c��O��;���~�#C* ��|�O��-|l����vWi-�gkb�6��e���~�(G�$��Z��e�t��yg�}OB�� =LВ,[Fy��c�	k�W�2�b�[P*W�C�z >=�'��ܩ�`6�ap	跘;�]�2�LH���D���IE�%����Ղ�^��i��f��F<����V��Tz���\�Ա�l�5T�)Y��lp�6�2Ǡ��Y�F#�^CzT���V/��.�[.�:�n�X?A�\�4�!�=��]NRb�l����z�!}$�:t�-%�U͛�7��&�z���"߼+�cok�F��/[�i��7Np�2x_��d%�!�z�ȥ%��x��wd����d��a��"b�2&O��d#kG|5���A;��<�'9���D�6%�l��Zf���*��{�RO9u�Vt��@_s��X��+�n�WA��r�_u>Z+&)^;C�� �=}�y1���53b
uՃᥬ(ߙ�����/�����0!b������Dpq�/Ky��৸�K<l�]�>���h�9(��Wg��|@����j��/�LL��⼂����\��`Y��:��yE��N���>7�<�X���q������k�n��5�Q���$�Jrh�)NL3ٜ�����T#i�E�?��!�v`�.��f�n3?�����d(R����1�p�*נ/���!'���F�����+8�P�la����~�w�n쯫QJ�0�٨�t`W�:�k��]t����_��j&���uQuO��+(�Bt륆Z|�?�]��`o�Ox�~n��X�ڳ��:ׄ��q���In���
H�S"�����4�G��m]�pֹD$O�N��k��UC�O�@��X51.�y._��&"!�Z;���ҍ�(���x��G(���̾O��T�ͨ��[ݶ��c��P-��|u�p������J(-�a.N��Q���2[R��u�j�A��О�H�{f���<ͦ�q�oyt��ɂ�O�ϹL�����rJ�(���>���{���k��Y�f8I��!�e�& ���_W�W����sq�k�Dv�GFq�]�Τ	�v_����noU��ʓlS��Z�fG��A@�mĳ��C)z�$�w{&@�����ju�u�Ѣ�4���]�-�����Y"��(W
��~F�h���>��#��e�m���vKɥ�A��5�$XK`B:�p�ɖ��
�^9G�e'!ۙA���Ї9�	���+�rNA抾�⫂��WT�gŝ�9`�b����X#�iq2O�\Zv�B�3��@y��k�FO�#WT���� 0 4fsT�TK�^^G�F?���A ����J��_�#��x��L(W vY6�;�&2Pt�'��=��Y.���G��� ��I����Q��w��|ט�~d�B�B��?���͹�=s�Y!�S����s�f��f��&�
�4�J��]�I�[<�x�!9�g�>�I0����hp6�,s��ȼ/K�
�m�Ie#�S؋�U\X/
�#t�ڴ7� �1u*�}Y�k�t�ܓ�'`����\I�^��Yҗ�����4�<�}g���b��>y��`-å��ֺ��?q�~"�-��y��H�$>nˡ{�-�ѽO�P��$hz���3���0t^���ļ)>��&�bm0�/�|ж�����.Ƀd�D�� ���[m���L�5�Ixn���QF�"�ASq��fs�H�(ܚ�=׾9���ѕ���g��˯8g��"ݯc��l��p�
nn����騐��L���X�Fu�P�{�F��H뙺!��N*P�h���s�+x��[�{^�Z���S�MNǁ�H,� �MQ&��X��^��6���������l򩨝b��ήE/�wr�0�Jw��}H���OQkb|��T�m��%؟�y_H�XC��_��A��'�����G{^�_�����.A���,7�ôӷ��Ƶ��ѫĺJ�%������XC����V��g��l�l /I�2=��<�	��� ��.V�[|�c!�8���8�U1�:~5D^�k��R�l"��i���^��&����̳o>�lǤ�d��bT��X�o��P�]��?Aq��U���)�ޔL�Ə����lZ���$�A&������M�����r�'�x�>�$��8s
B ��f'�fS�:f������͔ڗk1�\���=tSsUP!�W!?�3| �);��6�@#8����#���C��'&8O���:��Up��q�����IЙ�ͅ��W��+��bh	����T,��Ue��v��E�mT�����-	3)�m&�& �׉�,��ګ�c�����,󍛜T�r��&�CH�-����
��*�h^9���ل~xxF�����?w��S��R�r�)ޅ��)��lU�)�N�z`>�?W?$)A�F=�s�7������y���-s��N�ƣ�)K���U�܁C�4�jhÊ_��٘�h�;>̎5���p�Ů�O���� ���1(���}�Ӭ���ٱ�۲;�K۱�w�	gU���}Fg�Z}]����1C l�\��?͌Z9y34��>*a�l���?�8-f�s߆Ą;/��E��1��)m��qZ��M*dҫN�I-�2��$�)�Y+��� ����3C�f�H��7�u�66b'�ۦsnyL���:��#�[�}�ʋ�Q��<���QӚ@S�%���b����O��W{P��r ��
�5�����5��͸E���χ�`�ة-z�#�u] n|��Mz؝r�0��iy��w�)�����B	�s���V��*��9壜]� 8hFz��Bg��b(}j|u�b��5�����E�+nsw�*Q2�;>����Y�Y�����0>W4�v`JC��L?���b��4$�$ˇ�n�#]_Hƒ5�"[���&�`p㸅(���y(�k_?��k�T5j,��-�9.���F��O�� كC�$�%����g�rI��rT��ed�"���9��-�Q�~#Q�8=�A*h�ܽ��5}��eܶ|�*
Y<��v� ���e&�6ǯ�}���+���Yx$ݾ�/�PKȽґ�O�	��뻰���T
�L�"x{OM���9��,�_��L{X�POP�H�ywvR,Of_e� E�)"&tyN��Z������:���_�n>Ϗ�SY
�@$y_�PH���A9�3t�I4b�*zd!Oo�v_�u&s�٨���b�^63*b��HIYZ�w����s�OnC��{j�vF5y��꽖
���U�x�<�'~Ѣn8fp�Fd�DT<��j$���قL?�N��Kn�"���62�M �
qbZEQ�9?�.���Y��1����h��Z�X�ł���5�{mCվ{��	e����r�$��ⴙ�B3ѫ..ܳ�Tj�/2%b���e$���O�.t����� S�n�T�iwj��ݼZ	��|8�y�sF6���~��}�riU��N��T�&������k*�	���I�i�"�λiJYa��E��Ex� ��z�CT��/��n��Ru�lنa$������S��Q׻U7�N�E���[*h����o��ؼ �z.?��숢���#��bϸ~R�~?:����J��P�5Լu�X�Xz��)kڸ����a>�Nus-1?/��Nߩ��[]��.�G�4a�5��oi9�?���y(���ܚ�hJ�����Q�hy�7P��6�ڐN(��~��T��Sj~�M=����~�����od�O���d(�0���_����"� �h����8l�겷�=����a 7?���6l��i���?��	�?X��r4܏p�_���R`U��i�t��`�GF0�Q !(0N�������� _;_D���_%��[���4�B6�h���v�F3>f�3�lЏ&���	�M��l����Y�ێ���z9T7����T�责�e��+�mWM)�X��̓��}�4|}���tq� ����m�&����*�I,�`k���QA{&ķ���؋�';�,%��
31ݶ*���<'�?�����Ȭ�B���(椬:]�0���F�����V��l�L��҇5�k���V��Ѣ����vc�u�r�g¼.g����u�q�ݳ�VA�jf�}���ʁ1����	�10�K�r]��W���8�;�i�����g|s�'8o�81��+�A�B����Ω��u�<ay���������+B�1(h��Fk�u�\)۱��o,灓ԋ��PL�c�:	�����;��n�����YNų�=T�tV����f��{�<Wcr�)�ɔކ������"- �|Yb+	�|Rz(T�S�/*n^�U�}��E��.~"�-��߯�RC�-��V^���,:�>�S�|zZ`O��N1�%X���m���6�>�~}�(T"`���h6���	F��h��,<H��5��Gq(Bb�0!Q�2�D$�w}� ͖; YS�!x~����F 0�6�H�*3�h9�y��_�W�ʟ���(�Z�wؗ�C�Yn����W=߇�����lo��r5Ӯ��f���Q.�/�p�G��tk���"�'���r]h36O��QG�$a��:${�~q�m�1/	و�� =�������FPD�zXc8�3��yy������~���)�ư����}(��J�t9�/t�,7�赁�s�����c��?��b��7�qs��v�.�'�wv(f $P*n��J�b�����"��#�ɥB�Z��h2����S��_w�� ky7ǳ��JK$�������Ϝ4�&;W�X:���ŀ�\��TY�����-��89Ǭ�Q��N�P{ '�s�v��ձ�ty?3
��	o�,���C��ܯ�/4�R	�g�5�}k���s��r��<��=k��g� �mAh^�
wz�B�����������T����C��x�>!:J]f��]��N.�`����2��b��T�"�s�$\���ʮjLF����򒥥�w�d��ӤRjT��J�a�-��-�2�pA��T2{y�?�l,9Kp�#����:�(��ޟ�߀���_$��x7����cmE>����[f	�/U��T*�ٲ/	�jq�5ɱ7ϼ�4�&u�1W6���v?Z;F�G����kW�e�$�rM%����^{�l� f`��I��l�}z*�I�£/Nt���E��F'�,�X*���`D���Dхh�l�r��x�0)�T�.Ȥx�8�c�	�����x� ���o�\{Ru��	����@���>W�̎�T���:�g�!~���]�|��m�w��<cv}�BVw��\�u�9��lnce&����{�/T��B"Z,_p�gro�ɞ]ֶ*Ίd%��y�g[�����w�E���_�����'���d�NH�YRR�[��Y<�%�v�>�2�����I�AA~*�F=L�B�m��F=�뵍��>�1�P�\m0�UG-O���u���J����&j�'k�m3�.�3B$���x���b~���3���tJ���{���`ȓZæ�F�+���ǹT���\�QOs$����2��7剄e�!�i�xi/G۱�*���!0�'���D�̝��c�΃	o�����o�\]��I)���p ��5���:�D���\Zkܤ������}��Z��N�b�Z_�1�t*��R0�6e�"�&V��H_��Jwڭ.ۄ���%�[f/��j��R!���چ�c�|:��?nv@��Fm�N4#õ|(n�)x�mH֍�B�o�xn���#����eV��x��
��D�����������c��{�?�U�p�C�+Z4�|�?0qi��#�Fijka��"`�BG���9�YU��`>�T��e��{����>F�Ǫm�X�V^v!l��_�Nv�η�	���5�/�4�;5���M���N���f������|���ǢAx���K.T����*7����r.멏��SYe ��ߢ=�-w���OK��3��E43)~��C�!Z�Z(`_'�ZZ'g-���� q2�䉣�q}�5��-�!���9��R8�6/n��"��"{�b����v�S�U'-y�D��t@��4���	2���K$�\d�*1���+��*�G%�T�#��`�9�3�*��N�Ƙ®M_B�3��	�����O�J��w�*��E�"8H�+u>u���#����E���fl
w_�K��� ��ӯ7;7G�w�l��#'��3�5k�_L����3=o����!T/��À73��(�\p�V(��#�slWu7D'��`���} �}�?-%�;�_՝Z��Q���\��	��vF��p�!���WE��9�Ni	#�ǈ�/��\hR���;^��W���wV��[��������U�s�m�����8P�^�Q_)R��n�K��v��.����|��S�wK��1��wq���̑)ds��C��H���d�q^9�P��f?�_2�p���#��`�CY�q�fk(���ѿ��HȦz�%�u�d���(��(�����|K`��
Ð�,���LN�x�>�l��ٛH~]���b�[7��~_�=���^V�85&��C6xk�De�&Ù�D�R'c�� ��p���OmO�#��s�'�"��m�;6k�U<�AC?+�Iu�ˠ���ߡ��U�<�Cp��Y��7^Mȣ�`U�snk��a��;�R�4P� p'#������������*-2��^�j��ʀ�:S
��)�q�BY_�bm�&��^]�)�J�F��υ<C�/��Hb�>-�Wm��
���b2�@�}�m����ʘ�g���ŨƬ�6�����G�,t��=�Vp�(��%?��$�D4�]s���2P�G�q"-�1
 /�{�[���������E���J�%�r47�2y��!p�\�n����/��^Z��3k�Q��]����=2����[g��F�:D��߮K��������z�����od$�h��Jh/#A�q���:V�TpQ�u�� H'��h.��Z-
U��L�Sh������x���ΘDk�1�/���s��t`�l�8�Y��>:y�6�u�l�[K��3y�+�P����a�Y1��������������hS8B�2F����<\o'ǥ ���r��{޶/A�+q��>�<������;��`�'�­��Y�]/�B�]��Z�a,ɽ8=��g��D
�^##���/HW�Ȋ� �;y�	��p����%}�a��c�TpQ�������-��Y�>�[
5j\��� ;�F��6�r�HQ�zd�ǿ��o��쫎%�,���!5u��M�9�)s󛡲r��]��P��RcV|w�Ѓ.U�����oQ�!�;Wzo%V�����
�M�����sH��gt��Mx)G0��d�l�!Ĵ@E��K�^������QA���H��s!T���8�fY���^�� ����9A���n_ї��5�M/?l�&�x�_�Y���;�6.�Q�\���8*^P%�M5��N��L�� R������ZB� e-=�ܳ�f=p;5��d����y������N�Sx�<ڕ�/�V��VC�yNi`r�s����x�k�X��Q���<g�F� ��7�L�Ѧ��}��>��24͆+�S�yزx�N˃ÿ�kl�>�?v�Z�	�ts��)v�$=��z�vky���
6�r�n!���"������O�\�A�����A�-�5N���rAW�,m�%�ĘZ}V2]=�����w�R�>$���d� =]Wͼ;�uf��i���]��ZEQ��gTk8���w�n��0q�Aɉ�|�Y�j�g7��!|I���d����?,3�$C1'����I�L�:��-s�=�Y�g\��8릙����I����g�w��n��> @��l��;���O��9�T;C��ؠ(�Y.�!�A�~�@�8������Q��+�Dr�
�=,5 2��`Ё��ߏ}B��䅫��u�Cð�s �=�CJ9[����E�DR�"���7�����t	�e��I�Yh��\�����HF٪�wA#%b�t-�/=��!��Ř�\	>�T��O��.`HGv�H�������w}>k`F�>�����lr�U.�($��&�ּ��ohmL{}N�d��pt>?��̄�:0���������9��v��uv+��HUt^����;Ƨ^E=��6V*�RY�D�g��.|W)�Dl��$�T����xf�LR��<qxq�kZo�{���@�8�h�����w�`�v�3�/�T)�nD�@��Nł��2q]�}��m��nǈV�zXD��1c��w��$VA/j8f�� ߍo?�\َ�{a�G�Y�j`]V�r�2-��%�ˀ0W=T�* �U��r�&�� ��Tq��A��<�!5>��M��
`U���H������m�
�P+j�|"��YNO��`�Uތ	��'O0�V����v�6��6�E�,\ѷ5?� �a�R`�U�:�\�0��]��l՛��
؊�t�U����d^�+[�Ԕ\����UC7'<�&fݍ�!/g�Hh��6�&;)y'0҇w<�#�	�+���
��=�)�3���C.g��N�:��Fw��2k�!Q�3�Ga���O��J�Vm�t���l�ւ����8bU�"�.ɘ�V�FV��oD���`ǦЈ���37dBO+�E����IRԘ�*�a%6u��u�g����u�H�cΠ}<Y�����5$�/K�4��W˧=�����&ې����lpz_�����ut&r�%�wA��L�d[��^	g�l��_�ᤳ���G'��Q${\�_�����N�_Y�D|*��A��B�Oꗶܴ�����u�{��bV6$zL  ]��	�����"���-n��:`8^`v�doO)@@n�bO�)F�����\\�(��_`��gr'k�s/�S��K?-��$6E�c[�Z#�d��Ӷ�Q�jSD�x,�֖���N�9u���0NK�ſkd% qm>D�I������s�BM� T�y��*�qu�:�UzM|�	�i��)���E��[N���d�G � ?N��G�Gk��p�B��-Y�&3�1O��XĆC]C2bWg�е�f��0;��k6�Uν�)iF؍�u�j. 5�8�u*����RW?{����{hh1AS;���YX���z=�(0�[��z�&�['�tof��)�Iy��F"Y�������"�������Iq��:Q�%�sx��w����И�vLl>߈�r�X�Ug;l)l�g!�]z�h���|�g�>B��1���������k6��ʧ��s��?����X~KX��x�2���޲܀�;��b��>B+�cTx%��Ar7���[�T��H��yr���BL�Ӫ��5�t�M&�T��n.bf���J�5���fX�"b`�/�$�S�X~�]D�����T�׮��Y���{�m���/	v1E�gup::�R[L< h$"y}%� ˻��z���G�X�`	}�s���߃�Auk��sak$��	Ű%��2���v>�
��Q{2,Qd<-���a���$ %��A����+S͵8�݄�95�D{���=��x���Xy�Ϸ�� �A���"��������/��dO�^N$�'(�4V�/wx8��\��;^�N��[u������c UV���3&:mr��v�4}�t��o�r�xW�VLq���;	ϸ�K�����{oH��C�:�x�<�|��Õ���"^�+?I�s�0!��hѿZW�r�@c|�}$s����KͿ� ��B<b�1o@�/�2#)�J(���O�j,"�z3�h�Ub-Mm���1Ҩ��U���"�m��_bOr��BqJ����5?~�7����X���g,7�6o=D0RCb��\]���#%l��L��e�v*4���YI���Lf5��d>� ������I����4%��\�A�[rb<f��$�U͡+��K�A�v��6��ퟸ�	Sn�&�J�B���1z�H�;jr���PLzj̎+�Bsw���g�wۖ93��ۈ��cL�8�Iĺ��&�U��"�j*�մM�ğ��!��vSK[��x.�as]2���1�k�Z1��u.���./	Np�u|�RS6'
��X[�?:��~�E.1>�{���oq~:I�ϫ$����VgJ��h�p���Dn���ǵ0��pet�8�뜦$nE�����9�b�r7T�촩��D���7<�-��D�BRz�����Tށ��ISy�u��h�(���IH���yB��*/]%�
�����㣑q7_��>H˄������K��	s;�����}ޣ�@k�S�ô|w�1�� �{� T��mV������;��0��x��.3��r��/�l۪���w\�2��D��>~]�)1]хS��EF���2iM$J�T⿲�{ ��%���_m����ɻ	��҂ Q��hPo�d4��TV	Y���G	��4/��@u�k�I��4��`gF�ˬX�Aqi�5�p��Ađ��ߑ	�[�p�Zd����TT.A���V%96�����S���Fhx�t����=N�f��Q	��y��7�ȟxc�s��t��W֔>&̃�ŷ�)b��Fۋz�(��<޶��]�J�*C�=����d�����ߣٚ�S�
�"
>�&E�#��p䝅����`w�C!Ѹ����ՠs{���A
�f6�L�m�';���CF'�X_MOԕ����j��� ����$�5��Z1�jk69��^������}Q�q��z˧����t�d��(Y�{<u��wa�F��vt!�r:�S`���n������C�A&3S��
�L^�ݓ�.%.Ԉ1���a9��O��M�i�@�v���M;H1�]��h�bev��ѽe�o'B�Y��f�O�fr�e�A�+O��J��޶�t`V�d9�o�._C��i{�ΤZm��!$Rv/D�ܛ�|x�-i�bS�X82g"����d�,�?ZucO��~��+V	�sڋ�#�{�s^����"]�%�#���]�l�}c� ﷉����D�E_Nr����?��9f��K�H��2�%�;�&�O��h�l�����^4۬h�z�L#m�8lC��]�b�˹{���Z���v�U�- �ò8�R�6����@��ܗ�
%���9p+qpJ���M��?Yo��p�JP��ҋ�E�L�9�I����hSlU��$�(C1X�.��C�H"0�C���7F��{�����"(��V.α[G�1i�<���4������ڟ\ϗ�H�D`	E�C�^��h3��ZA<�ܝ����>� �D�ʄA�Qز��Zk� ~�RDζ�
2�V���T��2�М�ú��E��h��se��G���D��:T�o�'ƶ�����I�.�;R-RoJ�˾&�i���Ƣ[p$VK��#&!Z��%�[(�����w���,�:w'W�����X�I�%ۨ�O��1�����-�P�Ǟ�T���04��9���J�a�]�{�	�9=�j�ڬ��Dj��ǟ�Ѓ�k$�v���{����G�-;��ê�����S�4m
w<�ï�y�~�!-�ߋؙh)��J�<��I��E����w�D�RXs&����lZ�8�T�!v7�޼���X���r)L.���~��p�7���5����75A�o�����Tأ�S��a�	������U�U�D@{�:�������2U�t�$e@oD���oQ"�xF��#�@�����А���pYP�P�1��>��}L� ���P?�����u(���l5��H�*��d�\^!.���,$M�N��6�T�C���D�o�s�Œ5D��6#�`�|ӒT���f�v9^p��5��Q0X7���!�~`������l�Cs ��g��>z2��T�F�"��;�
�Z��p;iA�˦.b���TRP���\�.E���_�w]���Ťe���j��i�]�3Ц�d�F����Tۺ���(�&��`�{�2�v�����^��tn�	�Jq(׈�P֯��r���M�q)�[爋�a4	
��r�52^�bf�f4�o��	�k��s#�������
���_�M��0���sd�A;�w/���+���=��U�N�pqS�T��[6u��iM%�bƏ�M�����+��Df��n�D3���o��|����W�dm/߂Z�]�|Kmla��S���.ˠ)O���Q���"�m�_�/a�/T5=;/�� y/o�r�ʢ�lW�QH=�ӵV`R�q����FH��~�8�@�� ^��P0�j�)9-��k �����׈�Kڟ@ob���g����lZ1�Cv8�p��p�b�L��郒�:�hT��)��7�6�*��asN� )��U��ɖY`�E�L�F��_!���4�q�π>hB��V�t^>d/[��.{ ��gaM)RH�G��h��V��ᡠ���^^�h��ɧL�M�wfS.�7a渔��P��U����q�Q��%�����9y��k݊
[0�D_������ϴ7x��x���2���'7����Q�!�����Y��f�з�=�P��,޼;�(�a���UFh�.l�ؚ��(�a#�V��+��!��;��Ģ��l�/�̴K�ɗ�\��p@�	��g��D�<�3�#�j�mj�fy����I:��5��q��Iq�T�] CB��a��������mJ��U�9��d����kz�Pk��o���jU}i/�Gp��׎q�Pȩ�3��w}������E��^��ū��1t��Y�~��]�����ֶ!��U�^�׏�����(|�Ua�t}�.��z��`��no,֔��-��S�&\H(���[���-�2T/��X��beT�Z���GAvd>7�GԼl9/Q���yj���Q�m~�C�]�'?���xZ&S��u@َ�^��HڞZ_����
2�|�2��������p��� �Y2��� 6����۟�l }ś�R��౷Q^��'ڋ������Z_.d�Se���F��*G�M!x���=�I?R;�^�W��؉X�I���'֣�e	�#�S4���" �E{hk1��>ÌZ���nx�6u�T��i��>/;�c�@�Ī���bg!�6����3�|�Mtw�F��]`\�X�M"�+˰
�� �1����K��w\�- ���Wb���Xv���}xbQ�ru��`�@C�<œ�$G��p�N?@!7
�w�>��h����\�_��k<D!qS�����X�b6��{1�ur[:��8��';��Տ~�ɼX����[q���L��	�5���e����e�L����]zSc�X�e�>f�C���N+�ÝJ���n�&��2+���3��N�J|LS_��pHC�
"E�b�sH�27�}tg��"`�L0ĉ:�9"9z�
I���DҀ���8	�3�����wj��*��I%���L����if�ހ�t @�o�@��7�<��z��d.j�Jf�oP��መ�̏r4K�0KW^�2��y��`�5�ei._��yʵ���@Vj��oX���{0�R���x���m��yO^�?�)KG�ⶋ��ig�R�a^�� �r��@�> �� �揠�t�w�����\^�K������)�rG� ۧdy�A�&�tOh,��^l���{ALF#�laCO=]�ڸ���=Ĕ��� ���Z�ڄ�jw��(E1�/U���dYr��	�ڨ}���	L�a�a����kއ*� `W-m��;��\=����k���1|1n������h�g�ʛ�
 ��;5��~�irb�d����{�x�"0ƨ~n$�B}lv؅���]����Lh=�γD��9����	ct�I
�M����V��z���"8�Bu�<=��f�zH��u�6��Iom��Z�B2�t�ц�/�ޱA�%�� � �5��oc�����޻�Ԓ�8��(�=cuZ�`�j`�6 Z\�G�����bS6��;����>��yJK�Mu�H���C8�l�ucMRP���D!OSިF�&�>k����=��Wc�.�˄v������|udI%���-W\�Mĺ:�Pp� �l1�r����c�Ы@�NR�Cϐ��Y�3E`��_��_�X���%�����gSZ��G� be�����I�;߳=�>α� 5�?7����)v��e��CLF�����iλ��8[@4��	�G}�Dg9GF�ܹ�g�D`sk�5-we���-R�K��f�F�%(�>�һ��+	նw�^�˺n/���h����4�֩���1k�V8"{����{��͙�9��~P|Ve��Q^�6�h�ȸ���u�R8cՎ��[%�j.	r������7��R>	"�o���/��@��t��ܕ������2w����6��i�9�����M��]�ۜ E�i��ap��}.?�z��[\?j}��T���?��-�m�C=��0�)���%�.��R���dEBt�e�&�\�K��$L�S�i}�E<�˿�{4�.=o|zI�_EB�{�Kғ�I��gpI��נ���ɔ�<`�ҥT�ܪm2o>h��U��I��}�A_�p]|�d��� o�J�)@���c�{��������Kj+i\���qmܲM� �J����p+��$�;)gП��MW~�Bs��7�R��9��K��=�'� �N4�Z�&��=�~����g��a�p���[M�
���~�X�@V�����$(���O݉*BE8���\M$�gm9��Ү���(��@a滦�������t�H��麅�2�5��+�{^�����k�Bז��{]U��A�z�.1�x�]�s���}���"F�`T���O��ӝk�$��3�u�	�U���Y�d�B�%!3pvDj@�&��P�iH�������@��Ϗ�&�1q��L��/�k����V<Ԛ�#͚jl�?}<�t��.߆���ˢĔO����զ�%Ό�m�
.��,<���o!K��]=T��$�>����{����6�P\:r��sq�}�c����+�B1�I�B��5��8��w�f"{5�	�|���)�@�n����t�m%�Y�VZ0�c�1�Kt:� �9��Ǒ��2����7��-�lډ�u(;#E�gP,���c3ۦ]7�X2�7���{�Y@�k��{�b~�<\�z����D	{ʎN�K�+'�⏧�Cq˻�;d�%+0gՕ��-�#d �͟0���v�n.�҉�� �B��	�Z��
�N�y	.و<�h��j����A��"d��L�_4Rʭ$T���5��wf������w$�߆��{��O&,�]�oi�>~w��HU2��]�;��9��2���<'\rm�Q�Si�"Y��70�(�����yurZ������eP)����7��f���l��Q]ρSa�e)��7�F�j��`�u!j,�BW���
Q8oJ��Z,.���4�R�������cX>�3�8��5aZ~3[�"'s�O)y�ԝ�{�O�л�0(¼��Q�32��S�-c�m">�C��/\-�E�L��p�9_�5�����1J�L�-��_�͎�����VB�������>gv���.p9U����Z�_����p{Tr�DZ��i�swo�x�I���T�ѐ9��+��{`&�A����mM�F���qs
t������>�fّ��.FS�� ��E+�w�~�f�c���'$)7���s�5&\���AQPĠm�3fI�Åx�~m�H;N��\ĦEp��su��F���j5c���$%38��2����^$E~	&�$K�D�3 HR��~ac+#�x�434��� �����AO=�&;�M�H-\�O�ݥ�v-���*S�0B?O��w�W=Ld/_����S��"��$̤����s+�_����]��!܃�^z+~1/+E��-���L����hK�j�n�GGf��I���A���=~�+��JP��+G�U�a}w-!ѵ�/�i�\`�<��؏D�(��O�vL>���-�Eca���w�ܓ��G#XU`;F���`]�����(�
�r���� �@��\.2-r����fW��<ډ,1V�.3<����%N�Q�P_"����Z�G}#���u�\�dU�A	���Q�]Q�����N�,��q��Nd�`;�v�|�����}��09G~��ݲC'k�dTȸ���8;�َ����L��	�d�vZ@/��-�t3b��D�)����������҄�-f��4�uN6A��Lr/�7r;��驾\���0�A�DI�g�w�sM�p1)c<��A��{��\ZvV��%T&ײw��މl�L3�	�����*��&iaȥ���E�+�"�K�HN2�*�B�Ҡ8�O�����ȋ��5{������ �9U��
v)'?wl~/�k:�]�pY��z�>�s�;IX9���J�m���}�/i�r��c�V@��q��sg_  ���sX������e<b�*l�x�#2Y���(15�!HK߫��up��}�(F��VJ���.m��%9Z�HTL�Dr4@Ji�zC��.L�~��p#��y^'���ˑn�R��m�^(Uj��}��bL�����z8/f�mw�C2��־� ���"��NR��p>1 ��}�c�vk���Xa�*�ԝH��!���;�&���:9�K۾�Ņ�k�~1�\�<���t�r�s�#��h�Q~(>�!B*�nģעr�gCk�
,�w�	-z񳫟S����ٔ��$e�;/�F�BH�r�������-�l�M���<�ɒK*��?J�eaB>�Vt^�|��h?�\�uI��WA��̥)�o� nߦSlqG��+-���M���[�@�e��(���'&��'�����n���G����Ȕ&�H��O&�b�J7̠�ʞ�l@~�	�{�uSo����ԩDI�_q���!�a���al�1G�q؄��A�X4͸ɝ�G��0u}�c}�c}j��:�=�[
z�?3f��{%��P%]�:��v�e��nJ��範�-��=�cO5JG]�~�{���M3F(	��Q���������D�2�%�N�ӣvu3؀5�$D=�#ڨA�b楌D�&���:DG�[��sٖaצJ,T�Bd�?�x4���m��]�K�߂�ȭ]/Kij�׌�ڶ��{�(Yj$K�+��W�X�`2��1���KHAD_x�%v�d0'Τ�aHU���O\�( z9 �Q":���[��E��=GD����<���f�(��|^�p�X�-W��ٞ�YVw�W��j`��e��nƹ�1�ٴQ;� |��q��9=�D5�ɂ��KjQٖᑞ�>IDV�TY��S Ej�d$�ٖ���$�/Vg��DcC����F��D�gw?�x�}Pbܻ��-�ʷܥ?뉒V8'8Rs-M��u�W3�0�4P�*�ޝ��gz�/��(���V�d%ޱi�uU�q�wv�!�/r��N�.Zv},��R6u�x ���y���+/���ᶑ~ذ��P
�	��jg$(��2l5��Z���t�q�\�-��pT;������e����V������`�X^��CI�J0Ƀ�z�L٪@^$��̠)��w���1���,���x*�>�Rŝ���t�9���æ���O��E-JBD<̉
2�d'�{ߢQ@�x��Dps�� �CDŌ� uj텕1QAP?�
��u�=-�_��.[�?��x�db�IM�X^Xv/��!Z)����i{�lq�_bh�����7F�U����v���BS�U��om6'm-6�w�Fk�U3��b9�m-Y+�_�� TY)d����W���2O-'�/�� ��O����(h'7�4O.��f���1�B��p<Y4���@�x��#�_�m������^��P�2�*}�����m��L��Yۂ�Kb0�a�J��:Ҕg��W�[����&rL�_����;�k�R������o�{nJ�2�>sK~g�����\�b�vk*IO�)�Q#���|���V<�1�mtܲ}H�O[3ӳ�T��6�}�K�A'�>�]����0mFCg1��(��'�<2˩*�kV��cZ����������k����YXj(�w
�$�΃�)l���U���{�r��$�����8XM��Ђ��!��Dw�|OĖ�5(�P����K3�j}��ys����?�����?|k����9��N���	��X�ia3���U��y`-�D����4]�X�'��%���a�E�?F��FBr_i���%9�u�Lz`��K����L|l��/+sHu���C1,��!�b�Tr�ǂ���� lW)��:sƺ;�׆���b{D9�2��eSW9�
�i�7���o�p��
z��ZHb�T����/VN{1��� �6�Oj�����ӊ���KT�gCuD��N��0rm=�`���*||^��>��m"��qn�K��	4x�A�׶��ٳ�f�ؠ�I1Z�]�hY,а+yK����^S��,qF~��{~	�b̝A���S, F�'_ֆ/,��FM�#)����/7�#Ïi������b��i�6�uP�K-�{����{.F�H}c;�I���Sd�F��k^��
9�VWD(�2�3�xr��׊���H����`��SUr��v��� ]|��;s�a&�b��=�����H����D�r-���ݲ.:����p�Ƭ�f�D>��P��K�{��nsw��ڀf��pj.UTØd���%w�[����;J��7E%�eH���y��h�!�ٛW�i8']|)$�IUI�Ҡ0p���$���kYZe�Hp��hL�\	5q��n�ٲ1�a��5�tC�H-��2nd<���8�#��9wh&�y�۹.��Z���$�SZp�x�u���j� E8�x�����`��S$-��L$��'��E��!��sfNo�����GG�v׀�������=�� �>��;�X����g�h��|����#�>郛����A�V]��ŷt8�Vd��ǥ�e w���Nil��j]��jka·�[5{!�(�O��&,��ԛ���௔k�+;<|.@�$�H����!و �Ww1Y�$Z(�� �mz�W��/��Ǟ�_�Ev�eX�a�FF���<� �}�q�$�'@G҇9�gW]'�u$�l�h*�X��7-�jd�������uT�xc���aO�l�_��m��������y?�ȳg0�CL��Y��"`�[֪H�\I0[�n1�lT�M3����O>*�Qa�Ղ�BИ�� tG�+2�bF�~����I� ��f��%����c+I���2��Iu�ژQ�t�c@��c��08Y�@�&��[��b�
�D`������v����*D�LO�����Y(��awr�u���r�E^&�^���+ꠁ[�X�/�\�����?j�$��vopᅗ�Ri�W-#I��6�#�n�KxH�I��XPo�[(��T̖G��1Ġ<���x��D̹M� ]����&_c���H�9] �:Ҹ��Λ�F>h-�%m_�ک.�U�ވ�O�;� �[�&�q6/����؂WA_p�O �-�[1l�G/z�� "��'s_=��%�
�H��@��B�ƚ��X6x�T�2�~��So@I0����A\Z-O\�R=Vތ�߮{2�����7�s`��Չ�Ӈ��h��t�m;+tQ���f�,���d�UsYi58�W�E��0Ķȿ��UAK$BLh��rL�+m���ٺ�.��y̅'�����4��2�6Ϣ@d�δM��*J7� ��ʥ���wN�(�Mj&g��[s;٦�G�Ѱ-1���'�V��y�tx�LBS�J�(�^_����!���tUR�W	��� 'n��[:*��/:��#�z{>r6���r�ͺ��fQ�$Gʼ�L��4���.:a����(Wۯ�&ɜ�n���V��B�
�LkB��L^����WhSW_���˓�v�A��hy�¶��uR����!���L�9���ȱ����9�5zuvJ��C���$��\��%�P�?���˯z,��U$��";DO��1p���
���GwO�̖A��5���'�W� ����'�9����H��Z
��T9��E�+	�Ec?k��V֬L����0%U�(B�#���S׼��!���R/{� h~W�;��P�a4e�0��U����8�{��`��B%B�8�W��B�Y�|j�I��""��:�>GR�^�4E�t��V�n|�.8��0L�a݉�h�wE����
�_�����;o���9�d��돣^��x�9��p~^���9��MK���f!���K�P���9e�3c:�8�DZ���ܟq�t���N6�ܳ���-�}	8M��pfGjj����wn�ՉN���v�Ukj���#�$5\R�TeEu�2��U�#σ����;P. i�f�׆��gQ�6���G��ը��`@x��z\5 ˢ統P�$�] >��<�y�5U:}�mM����8e��[��HC"�Mm��.�d+�)��T]Qw���cI�`f�ߒ�z�E��o�S�U��;�Ѐ��.{2�5�'�����ݗ��D��@�?�r�fFx�G1�H$�w�#߲��f���r���`��".ϷR�p4x���x۶9����	���e+���hnb�I��-_� �� ��_�{����|5(�ꆂ���-L��"9�n##ѻ������F�PrzqԮ	�!BViw�WNjjvҌ���2g�����$�������?�Ih�C�]d���u}����Gg�.��m�P��R51��f��E7�$?1�����Tz���$p�)8|ݥՑ�å�@��=�5��h�ȧ���Y4xl �c|�F&�	�<���5�M�?��w�����C�r�l��rE[�R,�Vc�b���f�(B��.ne}ji�5��i�DK�{8���l/��5J�A�J������>̲,����
#��Io����E�x�t�~����qn.|!zI�����[M3`[��tS|�Oj
��[-e4��>j<�8v��%(/8ޯ��~��ٛ�/g? $,� ��z�Dv[��ꛄ��$����[a$�3q��t�n�r����g�~�D/�S�p��[�v��>��U��ĭ�a^�:|}�����WE��:
�F7lFKa즨_lG��,�V4�/{�!0m�VwM�Q9߽2��N�5>��_ַ�����'�	����p����!fL4i�M$�>|x�y��3<��{	sxQ�#���ь�,�p|�k$Ȯ%�V�!ykI�u���Kj���-6"l
���<m��u�I~�va���@���\n�rFź��.P��y[�F�@Vۺw�b .��N��!�H�h���Rr��p,��.I��JJ�;��5~6��/�Ƕ52��5ַ�c����7�G#Ȓ�\���B��1��|:�i�u�����Cy��N�٣T=�,/�h�c��M9�D��w�V_���`R�8�vU`(=��7�S�"zoU����8H@��r ���s^\-q{�T�	�����*r)v�H�v��~�c�(��Z��) 獾��,��p�ٶgMן�.��#�h]��T���]
�UX9
����4�C:22Ɓ��8�öj�� ��;��3C�(*p"�|�6����P�K��Ƕ/�Z.��-�PO5ĸ���8��g�O|�n1t�x���Y��$�qFu�b(o�<Ý�{��`�It��.���$�H�F����zJ#ٹ�m�6��:t�lKw�ҫ�	��4_��IV8���x��ƽ�CW��,�v�I�wu #��;�A��������8^I��R��Ӎ=^�͌^��T�8�&�(�Kբ{�o�2�$��6�\*���]��\�K����U��(dj��]���eaT�L���X�L�dFPh惤��1�.D,ܶ_���2�q�v�?\��<�*�ҷQ<�::���I���4c���i�U\=^aK۞�L� =2� ���V�=&��M�ꥡ�U������#��f�V�ϵ.��b�X��=����lf��=�e$-��4&��t�����Y�wt��R�X���ˀ�����X�kh���W8�/�Q�/��9���Α,襘�z�Cz��/�q��*ɝ�Wa|,M��P1�z���aY�̄N��z�8��sm�����^_8����6���-G6�7��4�z�v�q�.U=*�򔴎;�|Q����I���
Yp*fin(^�^,��®�rI�:��[���h�{R�M��>i��u�\.���H��5=5g@�������-k����E�F�낟N�ݻ���C�4�\����â���t�A�t�cC�ģB q��Dy%�'R���|�m0y������x���ܰ�8���ж㾑���ق�
���Z���dя��ݜ�/�j�8�	m�i�����;oG�:�N8�}�� ��/��p٨?���  4q�9my��!���L��� ����0*�����܊8_���휑 �>T�O
��#Y�s.G� b<�/Rlz\8��`�!*�nA���g�%��l@��h�d�A.PdePYg���`���? �Μ%�������fD����$�lB�Zf6�k�蛈��F�{*=�g<��Y��"7�����h���f�x}s�f��ϫ��Z�G���"����x�6�_$�zN�r�: ��j��2['��J�?8����tC9�Ⱦؓ�v]��)m�\z�כ��H"�z��Z�1�8��''�:aϙ��
1����mg�9ƴ�̄)T�{`_�r\�&he����Sy�����֗��o���QP0	P#����odл�޶�΍X��H�u�F��	�1b����E������l��d"wG
�Z�u'��Q�J'ϻ� [����U���MR��'gy]�_�3,V���r�Np�^�k�yR�"":B����>a���>w�d%=�	Q�Y8��|01i͐��fO�:�g��_X�NK�C��4;�����h�3�n��}�F����z��v.ߊDDoRtg��㥛�-��b	�w;F��5DF}�V�ﮟ��9�Yւc�*v���|��Dak��4��E�<�}JMh� ށ��|9�IA�9r�g^Z��ꞣ�nF+߂�y����.���1�$ܞ^]5L5"��-5�]���*U����A�G���uU��*vf"]�xޮ͓Զ:� t��Eяl!l-[,+�v~��$�s������6��a�碏������,'g*q�A���44�?��u�� b��~F���n=��Vd�eت��!���������/��s\m�8a�H����P�28Śk�!���|2,�H��V� [(���h��g<-��[�!DD��r��,8����7aC�j�?R�_m ~�����G��ٙ�Q��.֩�B��6ԥ���O�kE(T�\�<@v���Ou���w�wU���TMt'��Q�B
C ��TZFL��~��=�o�t�~�xK���lh�{W
��'#�TP���_.P���p�g����8%�Da�{��`t�br�h� �ꄛ��:���6#t�[-�Pu�����ԛ��W��*b�N�Y�dN<�)p���Pe�K,���%�IQ�u�e��K>`�ޅ�@�����J�'���f*z�Z�$��K��� h�2fdc(���/�As�A��b���`W��n����ن<nE�{%P���7&��0���'���ӡ"S8`�i�5�����+��j�J���~RA]ǐ������]��dٳL{�2f�}j����ĀU�Ӷ��\:�c!�c�}$ce��n4\MQӻ��]���^�ks+�7�G��B )��^>�t�t1)[y��U��ԍW{��]P�|9��#R+=�G������Nu�QB\�7���6��E��o���`�i��TnI�%���H�i({�&@��>c+�c�*>�]^-�2o�V�	��1y�B�իR_N�?uv���A��8���&%D����z^�?��R�wY�L.9El�d�i�!ӧ�F�p�1 Fc��F��O���W��.}q1�O�R��z��z<8Ϟ� x�F��v,��& ����ٶ&ؑ۶�M��W��v҉>@epYΉ�I7��20�C�0�p<WC��t̃�7�-��fl�Y!�-դ�>�{W4Q� �6o�U��w�`?��y3}I�A>�,�m�ߘ�)0�����b<�ȤM:�F��
�{������SZ�����M@����	��6��U�A0���N��xAFt oV*=-��>�b�+W��3�ֳڍ�N]�Z�Y��%l"��:�H�~�	(�q[��l�;�?�:$�
�|��VI'^WI7ͤ(�����T�����H|紾��(ӂ�E��-i tW`�q5$G8~J�ʹ�l�<����f�/f!���{:=�:](6 �72t�*������=�b@�O�4��]Ln�|p�k6�p��6�}�Nx`���R����g�C(�G�h���'ȟ����~��d-������9٨d��H���e F�Hh�wR�4����s�:�ˋ�3x��|���	��5���Ld��RaC[��u�Y`f��8b�7gi�[S�kj~��/���,F���f�*Q�� �G>Z�k�ހ?�4�α�������UN�H:��a1�}���Oo�� �c�rLC�f8�{5|���2a�^�Ço~�t�/��B���j\�����wp֧xA��!�fG�K���MQɿ�˵���M��..�=zX�VD�.��z�,/�i��4q��V�|Ҿ�xX��o�L�h����B#����#e��,��?$�U�}3�y��C�6�Jq�8�������������&L�_�6�Tl�O�<[/�Dj���v���k�+�,H���@�����	!k��Py��*94���,���GQ	#^��b��Ey�O"����`g���h�Ê�K\=�K��p�%�q#x�ܗ�H�=cgB�w��-Wp&F�Jh�����IHBP��)U?���
8`\j��I��o��-�t���EŨ�,�9@9�4���ޭ��N"�����a�6C=���q
��� �����JQY溗	Ut�!��h�^V�o+�ˢ���$��S��U��6; �k��y�pC��U�3�����z*��o@���������� GєU,�˶��ۅ
Z�&_�<s�=��Up�Ԟ��s���Q$�9u$J�w�@R!r�5N�qx I�(�!+w�zsW._l�+��tj@� W��;'@�U��̡��Df_؆Yʰ��_��~a�L��Q�a����=K�(��=�ZhE?�[���^F�y�]F�c��t�B.g��[8؛y��Æ�i�L
��4P
�qK6dԗ�Q1n����,���'@(���OBiբ˴�w$�6c �Ծ,3�.a�Z4J%L�br����2N��8'�l䐏�@1,]dκ��@���>����}����m�gA��u)b@`n��Z�M�M��ur%��Ro��5ܨ�ѭ�����=�ms.\�~e�{k�d�g�yjՅ�{���ŌS/���:9��#��%�<��Z��Ec�Vn�ƐjgXJM����s	׽��ES[B�|(���C���S�� ��05=��B|�����͟_�/פ����h"��5;fzl<F�\xQk_����':\h�Y`���tu�o�����-�m����c��b����Og� M���3�
�ɜ�u���M0�>��!a�j?@w8�Տ�!$ �`l�t��h�;�vI+��̸Q KyL��iLL�0���~�K�{�[阮��Z ��;�dX�% ��u�#6�{DfYs5Z�����H�Y�K1�bI�E/�F�3 ��iS���$�����-�Y�G�������+�,�.�/6��ݗ�6�����^�qHN��j$�1��Y�;O�J��P�X/�T�D��az�՜���������4²k�]"wM�W���%ǉ�
=��	�K{Rd^[�5�1z���?W�i�掕��]�ܴ��m̙x�n@+����'R�"����-�=Ru��� ��RC3.�r�򄌫́@�lf��L�:�8���"�g�"Jݻ�]���5O�#�+�s�;g��>?����XB��X��ǓV���������诖�"��Y��_�_�ϕ�66X{�{���~��cs�J&��l���K��� k��t��d�3ĆWKJ��;S1������cd��thuJ�܏��r�K>vջo��Y�&��k\�U�*�P��N�K�8�����ْ+\T��J����쒿��R�&SN�$���y�uC�g�����r_���g���/}�v�I��N�:e=n�o����|�EN�Ĳ���;F�#�O���KϹrR((�5��
��72��h�l���s�J�L/���/�~��6yq���C������ʖ,�)�;GQ��yD�J!�Xj�6H4P/�f"K�����F�ÿ4iw10;���ɪ����zm�.�仡��3�+A~q�şH�j��
�w��-���,7=�`DTa�1�䗆��\ei�&�k�J�8QFU2r����8]y��\B�1g�/���g���y�t�oL�$�w��Ӵo�3ʞ\�ei�v\5��F�G
�}�{�3�؊����E���v�X÷qA]y�����ߛ��1���>��δ'g�l�"��b�d[.[�p��[����?����X��B(Ι)�m���?7������F��3�ˇQ�[�>���X�#� ��hn��{�\�<�sI���Hom�$@�Ƈ�������%й:��e�}�k�jա̒�y��{\���o6H%��յ�z[�P�v�	♤i�]�P��Tzؑ�����oK�N�Nl�_U�|ů\sT�I���+
1�j�yLVN�KpJ���T��;���RA�t�}�l�GJr�&��Yؓ�[�wG�j�{}�3âOX ��BU@F�1���.�|��p!���ҧ�Df1�]�b�����Ѕ��m�&b�����2&�#X�r^����	��ϳ�IP��t֖aY�>A	KQv'C�H����C���{U(��t��R��_��7|Ԃ`V��.�xb����8��,�K���+!.%�P�l�`�a+��_8ˆ�o��C�'#��Ԫ>f�[L�{6�G��T�=�b�}9�i,u����޸:0�������.m|�z5���Kw�� �tr����G��U�u��Ov.����R���JўDV�Ƙ���DCd��1�-����f���`޼���(�[��8�w	n�zҬ$�xF�4��ee�薜H�W�,���ToX���W�8�,�߮+�������݋�l���v�Z���I��4H�2W������@%*F� ��
J�Z�7��ٟmV�g���?:<�.	�����u�?����LROd?��P�^�ud�0�޶�c�81%cH�U�ؑߖw��5��ֿ��<�����#�%�j����O[�R��:0����/wھk���Շ`9W,��VєWN�D�M���+����y��M�W2�ƷZ����K��s0�����
p��6?Ǒ��J�ߞ����|���J�@�M�����l��p�vL�fj���y���|��i��5v��H�Ze��� 3|���G%�ȫ�|�S��������Ċ��_V���w�	��t8��]�(qz��������vVy���4/�&�CmC���T��z����5�;��Ѻ���$&J��5||�Q�Q|˵Bv�ȑ�D�"=rD�)�)���~��~!L��3A���p���-�T<����@>a��R;�=���Ks���d��'�������gp�g��Z-�V��d��q (����O��M���x��Ҏr�SA����as�<���F��l��/�Rq��K����o����c*�?�:��7ί��*�VW���KI� �N�d"�x�6�ղ]%e�����,*�p��$8d�|K�[Hm�v�x1���alM󾟙<���z�>5�|W��j�
�b��`2�hάK�֓/������M�c(v��iz _������xX'�~Ճ}NU��!)j�.�&'��C̎9�YS{ǆdq%Ϯ�#y���	���1/P�R�$�U��@^P�g��,�L�&Bt���J5�Ȝ&I�uu�*.�f�3�=�l)�em8g�V3�s�׃)~���X�*�JD�sԩr��&�w9�0����P�$�R_9=f>��9�c�	���+jX�Y����2f񥏽a�7�(����Q4Mں�Df�, ��ь=��vL��u�L�~�I�:��(Xt\��{���\A��>S��AZ"��Td��7Sx:g�-oh��Rps��� ��ZU�y9��vĚ�r���P�`���k.	�F��Ƽc�L�Nv�����h�/+4m`V"�#��ե2�;�:�uP�����'q#;:��� ��D�ה��Z&Ҝe�s�"�hE�#���Ŕ�Ae���e�d����Ԟ%
�	@XA9k���� ��O!�������%h(Eb�U_��e��ubW����/Z�P2%	�nK^U��JY��"�a��xs��B�˔/x�a�?�H\m�maػ}��x�s��U�m��V��S'b��3<�$������ʏ�-42���G��Skm�c�
�����uk�����P�>v"�sn��3���?-.�u$�	���X��k��'t����ڡ4ft�`�L׎�.;+�y��7���s  b����E3�(�����(*����}2��yK\3�45�6����k��Xe����$8_` ������,!���*��#XQ;��,"aR��F�����n����D[zW眭�	є�g�����q����F��SQL���e*�1��29�c����r�W�q,����`���Q]]8!mӑ��M�T�A���@���z��Sqoe@�*١�QKIЃ����*�Hod�d q�Srq�ڪXQ�Wup�ZuyE����\́��fٛ���J�{�5�ux�;�Q�m�����`�^�Ǫ�X>U�m�Ә2蕿�ˁӛ@>���Y���X0{��8���I|7;Ib�����M	W��8[|�R:�+w�h��j�Lߌ{�`�/"�>������:~���]C�Zj���#V�X�{��$���g�;v�O�z�/MT��wO�'�Q��3`��,��1ʵ�c�*�a�}��Ml���<��ӕ�`/��_�S���OU�7���>��'4ơ�9S��nF't(���
Ͱ�P�tr��+�2�ιdQԹɡ�@��5�ޘ_e�Q��o�{	A�Pp��e,3��e�qI���y����(�� �o��4(��K�� �� ��EӢ>��9 �H�`�)*r�4���>[b�Q�N�=�A��J�xW�;�Vւ���}2��u�*�
�������2�	I�A����{[��pY���8��$�<�h&�����`X�o�%�[�l�]��:��k]�%1ap�h��렌6�<����p���\�D�*��]��1:���,:���J���p�5�����6�N��ąs%�*�K�Lö�N���p�b�n�t=4w��H=�q�*��l�)5+\X��lj�nM�r��/�aЧ���Gϒ��I�!��R`P�] �y��\�șÐ���%�/ow�yc\��a�Tm��eu���n������RŐ5�2���*y�6��,��J2��O��#���k=�i� @���>�6nǘ9"���:H��,r��_������Tϕ����9@wf¾�SpLo����@_�3E.q��n���dw�͔��< 6u.��֝�iZkV+`ۗ��������l<����ʴ�(7d/%@��v��:�-gT  k���U�\2BhU��y�(VH 5����$櫠��mFUK?ƀrv�,��C�{�n�Y�B  B����I�X��6��c�Vx�D����.�
7ý�8��E�E�&�et�ۥ>A�1d7[I��U.�Tg����#"wMN�~�?`v���v�Y���`)�)��Wu;J*h)϶�-�D%O9�)l��Д@]�oĂm�=��e����Ȉ's5��M4=؛9>�|�0 ��F9��0��]x�d�Oe;D�t����Vݽ��e�pV:�����W܉�
�׍SSA��J4��n�ҋ}��(�ݛ�z�%����ޮyQ���'��(��עi��y&��Cf�B�w�j���;E���2C3���"߅���}vsg�h@M �NsY�If�#λ)'8��:�2R*h{��Tk���>!)܎7���ʗi{��C�u���b���� ���d�����볧/l���$R�U���L%����Uh2�{��%���^�o�Ae�=*������*1�^�%�P�n���͛��N� �燂�E�E�)yPn i�&�s%ѽ���َ����x�M�V����nGИ�p�e�"�a���X���g6�q�E�O@�|r#zv���u8T��j&��4\U�7�|o����nj�ݴ,)�Pf�1w�Gfe�q$�Wc���+Yw2�+E\d#ΊI[3���R3��|�wpcX��=$>�$���> N�������!km�XQU8qiK���I����r��"����0�`$�{���l��jqD�3+�ʫ�鏟�Z>��v�	�a� ����"�����P�����&{��$�i�o)��c�4��(��O����v"�k�[2�K�R9��h|Ko��8�P�~�X�{?w#�!4�<�;9ur�b	��6�`#�q�����l� tW/9���~�5o ��ny��
=�#U}bto�IT��B��)"�`�U���~g���ʀ)ԁw��r�""�j�a��_�%<��'N%U�O�\��j��T��
UKgŁ],G��#�|JZ���6L��vOぴd͖�6�LU�CnG�ɰ+��6,2�!�P՗\[V� ����ARl;b���4�e-,�pm�Zᤗ́�K(u��	�C��xW�T3��c��R8���i�6O�Y?�#{a����P`<�íz���4��A�⤣H��вa��5��m;�t�j}1���}粃���7	B�O��{ƍb�����E�ln���'AvX�`t���p�9k�B��>�ߊ�&+t`��hg��#|�C,��v��ku��N�9vO8r6�l�ߠ`�lb���[�YY�@b����#��u���t�%��H��1� �@��Ŋ�,>
!�i�Lǒv��@Y���X����"6�~5A�1Q��X�L'%�aظ�s����<cˉ���$�ZN��U�d��[yy�����{��qg�g��<��=��A�n�����缵�ϖD��X�$��X��7P�Ms%g��"�A��C��Ϯ�S�wOf���@,)4jMU�d�ϚP^��s1���/2��x]	7������r��h��&�T�D/2�0e�b^��5��j��R�d������\w�QE�W��������^��`�V�p�V�A���;'o�;���� X?����A�m-��_���ͭ��.B���a��3���Pk�-r��p]�6U\�ĸK$����#5�Xy���I7
���yF'@;~�	��'��D�K�����@Yz�F��A��&�("=-�<���_(��>U<�#�c�����ER�/>��r(��i��Z>��0m@IP�gtI1Mi�N���K����Y��c�����'/���R�i� 4Nv�5�!+��d�!5[Yʘ�n��4�Bh� nA��8���W�׍�($�����L�0�c�%��m#J�,���P�bok"�r
)���r����u&����>�=���m�� ��Qm5".Bh�-�(e��F!�^�h_=x�Vs�@Q\x���))?�ޠ���z��쓢Ȯ��#��>�4>���e^�I�Ӵ����R���I?�b��F�բ�b}G>Cs��:۽t%��]�C~���f��F#P�[,�yz����qh8h�<�ۻ췃�m����T+��]^�\K���WiM��TnY�E��'�J"�_�<\p��V�$I��:M��-w��0�G��Af&t�+��E:�:���ᢓ�+P"�^�p�f���E��f�5zi0��^D�-� �3��r1SqO�P8�Qj��-�s���׭A�#�ٕN� ���16}wd0��d�}�2������H�/Z�û�.�ٮ!t��]�[ƫ*�#��Hˢ�X�s�NX2Մ�],^x�2qS��� k����� w�_�)��_#��^c�"�rkl���e>����48����~"Æ{�u���G��� ��U>����u�y[<�o��ә*
Ȭ��*�61�)zqF��ۊ�I�R%iy��o�ۊߚP��(xrO\W����`��Ÿ]��lr2�W�Z]��� ��^7>�L4囏c�9����4�R'��`�C?Հ���0��'�r��rO��y2cgm��1A~}���tNQh
C�.�BT'�v�H?�������i�ݳ��E�,����>�q���i9�-S%���ۊ|ܾ���T6�nv"��Cѹ��j(�k�ъN����bV�b�Ç�7cq�v�b`����.h���˪���&_�h`�~���a?�Ҫ�R�yx�s �N&������.��.k��t ������(>��u1!Ʌ韛�ɗ霌�ʜ@P��CФ�6=�"���f�h�nl��*�~0��|&*��E�>��ʊB��!j�0(YX� Z�� �XB�œl"����$!�+�����|g��ؖ�d������rm����r�r�V6�=9"�GG��Z$��_m8&�%�2�c��E���x��E��D/�-{����*������+�,��M4��ް�]���>�{�<��>3t[�A�f��0�D�X&�{�F!��$���ŝ��M��a���a����C6s����\�-tP�O'�p*.,?��o䙤5�϶�����>��3��Ӟ����%ⷘ����*�+r��@J�T��g�0�@v��;�7I\��V����<� ���0����]�����Jv���cq�$^/P��c���;��Q	���ON�~�&�B3`~�_4Z��*�*]]] �8�*��ɦ�E���ߌF�QK�kM�^L���Xc=/�ꘊ�x;h�[�:��{S=sP��[����-��L�9�@�������ceЖ��+�EӁ6a/{�e���9b�������)mu�e��YZ��6`�W^��U�����S-/Xf�ୱ�����sb���_�솻솂��rh�GW�0{>��I	��b�_qq.��N�c����d:��-�AY��]�q�4���D�6S���j�s5U��H2?�CxRY�UcX¸���_�B���~*/;�^-�Z�>������6��^�p��_�N�
	����Ul�5h�ڪ���.��(� ��.�qx��G�5,WY�n�e#��j��O6:�AŸ_C��M��c�pP��A���0�h]�s�`�`�
3�eW͎T��<Q�vI: m*|V�-��K�JNA�q��+;h�y���߭����a�TH{m��[�+����y|�d;z�""�r�F2�E������>A.ṃ�՟ο˨M�D~|�G�"���_ؽI�q�
"Z�'�^yVw�W�H�t��'����B�N�:cűv�{��Xb1�2 ��s�ZW��!f��D�g݀`�m��S�]�=׵_�����(�Kh�ժn�Nx|�}%���[$�l����9�t,���rk�=����\��ߠH)�i���X�&��T����RGY$z�d��, =?�	3%PuVU1Cj��$��з���Yk7�n����=U�d#�]�̂f RA`2�I��Zt��B�_��@���'�}R�U�1]�x��ߌl��2��>�]|5���etE��1CR�����z�[ă1�bI�pޝ��ߞ�"�z���4��{[�b�����������Ma���I�nh�)���~2>P�dx�>�/����E�j&���5|կ��@l���Fҳ�?Uo"/����F3F��I��ր���?��O�a[�U!r��_1�qL�M���������j��8���&$3&�[
���}?��(�)�Z�����Ÿ�pY�Q�'U�,�z*N{�o�D���rLF���3^�/h��&%P��m�aB��Ts$��.J��c(}�����x]?�ݍ1�sYե:~�WU0@g:U�lOM僒,��ԩ �?S	�Hj;ZU��n8�^{�M�$���+����C�`+Ow���,#�Mf�!��K�!l:��]s�
�a�������˰�.& �>�������+���Ka�J���azsA�k�g����[�a�pO!`IݪbR�|~�{m�P�h_'�QM8[Ca�3�����*�{��qk+ �H�����tvk5��7jɞږR2��u���$�J0��G�_�v�4Ʃ�m�>��^�:�@�bilJ�6;�4�٧q8��s�؆��@A�c������
�t��A��Q�}���H) ⧄��[C�d�k� ����X;CeI��9�Q���y�7�L�VR����ю9���}�����<+I�t��Ja�=n���٦�'��$PMV�/',����N���z�v�����5�i9>`@�\�o���l#k^]��X9��������'��uo����iiX0უ�8�����%�h2ڷDBx3��S��EY����"=:��,X����R�#��q�_i��4�3(W=�����D��$�G�LHΧ`��^���7aU:�?9n�,�7�o���d,~Bm;�΄�����
Em݁t�.a�'z�P�g}x�:#t�pyU+5X>�˷r"7��|YӁ�T��-5-1�5�~�Ҽ�0y�Ä2��������$q���?}�Jm�t���v뭧�e� P��vܡ�7ƿ@�ߐ���]{��!�Xt��-�cJl�[��	o|G��U��5�39�J}⭒�so��V�kH���{�,�3df�Zr��k���vu�y������a;a�ͯ+T�=���qh]��(��%aӔ��0����P�7�mء�+�/9��>�z����-�����x�\A����B2����Hx������� ����,'��/{��AjĊ@�~�׈ ��p::XQ-I�J�?m`��Ÿ�?ZHzI���_#���������,�v�+�\|��_�̦%�^�5��s��PeJOa�B�u�>C�^�/�|���ꥒȍa���Ej�؃3��"�q�( ҒP�rk��d��;�D�ACiO.P@��2X��C��>0�3�7�R�V^���;?��"�`�R��M8$"x�N�?�+���ɦ�.��"1݈�L�|�C>��@]i�9��?ĸ�8@��>tnX�hN�Ƣ_4xW�'�W۩�a��8���7R�;J�֝qB,R��0�Zm���C�M���2(V�1��V��i�
<�M��8\�)�:��XE
�D���M�����*�v_����a]�ҧL��E��{ �E�y/Ueł����z�D��^'?*��@ξ�"8*�xjD��)������D�6�:�FJ����| |	�������AVd�,t�B� L���rvW���~��r�2�/1G�`�;c#T8�.;B�H���z�:�j�$�6�j��v��Kj��-,��RÈ1�`\�%�RB��T;Q��q�lUh�C��GE�����ϳ��f���݂;m?������n�ޭ���R��a��~��>P֭�35#�e��@��ɃZ�A�֖`��|���3�C�邋Gv�U�:�A�P\����Ȗ�����-ia������ �F�R�)~�J`�,���=�^��h�uc��|����y?�}�GqI.�$D�_pX.��H�|�R7������ls�i<`i>�7o����S,����ڋEaxq����! �),�ْ�����51�H����v�ι>�tp�%A�0u�ڃ���{��{M��Ԋ�G�? Z����W痙���oB�
�GI��LG7�h��y��ϊ�5Tp�ڻDq�
A 9Yu��E9Ún����И�<�5ʤbp�O ���ߑ��+^_�i	=�&��b^���2 "��i�5��xf���7�r�Nዽ,#��N6o%��Xy�����I ��Wd弿򷅼\E%�	u}����)��a�|���{p�����C>m�>6�1
���l�"�!�?޿�.E��,"L����'��D���Կ�@l��
RNtld��p����\�s�`�j�K�����G��
�В2���5%Lk���z��O�|e���}�9&F��j����ֻT\�K�ѝ����4�a�%j���0��%}<Kt˗ �,Ci�@� T�1Y������D�F�i�c����Ą"�cP.N^k\8�$��@�r\+�f�y�$��X��������钥y߻�q�I�G�N4�!o�!�<Z��(�݊��^�&rG� tQ�n0���N�Wk�}�=E�y��G?�ު7�����9�ho�-5��~��I��>R `O��.2�5U��E�_�U(�G_��O�Nvg�{o�y���ѫ]�wӛ)��'x��;�����_��|pي��A�o�<�Q���(>,:kr��"�V���!�;�z�f�\eŨ���8(��T�	��:d�ؓ�~��u���$��Y,L��Ĵ�%u��'��_dF���8��+P�����īrH�暎�9$�9�`���wdMQZI�2/��"�_X2�e����l��af(����~�\�蓖\��@ۅM� ��i;�X\)pO6ggdQ8�� #.
n\Y]B�njn�.j7x>@Kd����ɫ7�YU�g��8^�%�C
���(�;E��?;W6ֵ"��_"���Y�>��`3ģ��3b���a��������"�(Bȝ�I�~��^�u�S�Gr��ﶩNW7`��)����s鐾�!zo�Y}�*x���˰��������@���UR�ٞ�ՄTe ����D�t@8�}e*�̩�J:bX��<�WE�~pqrU� 
�֥Q<P{�'e��>�gl1\_	��䅧wEt���.#�ZLI����L��_����LGhJ0e��MCf�^�ov�N�������t��_o��ONDߣM�< �'����4���E��h�I������Խ��г��ٝ,([Z�;r�āY��^*���{��}�pyz<����2��w���MvSrCes!쎴���ʚ8�&)��+A� ;
�֙�����|U��)�,��x57el�ņur1nɩvq� ��x ��mu���/�5�b;��:
^0�>�n��Bx��2��J\���ri���T�,���F��I����˙�H����8C���=^�1(J�G���7������ġ»I���32_���� S�{i�8���t��h�����R��
�
m�u�yϦ����7e�ke,���b�pa�w����gm��$�����O��.C6��/��W}ѩ��l\ܧ[���(1n�l6�<�%Rj�?�;�+�����ϒ�a��3d�f��%y�,5`����<��O]{�+&���_l�J;	+��@��1�G\mO��tl�*<��)��0{�^=���~N�u�`�Z������l~�|x6�ض9�ǘb˄��Nc���&�X��\��(����ڗ��9�8�T�}$��ro���:]�k|�oL�s;�k��P��H�6L;'��b����A�7 ��T�DM3�Q��Э���1`8(Ôf��ز�6����9K� T�=���]�}æ�{[C��-9;�I>�D�c8 "��̶;�����;v�3knZ���eGw�����b;[�����'��%Z��z��H��7o��M�
� Đ���RgD�-�K�X�D{�𵽦�h5�OB(<#�(���!6zjY��/�d�pQ>:\��KQ���2n���C�%F��m�d���O�����	N�Os�?�5Ͼ��
� v���#߳5]�:y����4����������bL��/�M�rv*�\+�R�M�s��#V���� ��$�Fg�f�X89�ԋ�7�@�0>e&ڕ k����Yy��$�Z�QMY�4�qf��(:�E�4��8�T���c��vl�o'���~C#���Aݜ���C:�C�a�>���_��B��>؛�T��F!o*�F2[�C��i-�>9���ɛ]=zR�"W�~���$�*�H5V���<�����̪jw4�cN�+�l麷d�E�F��-c���b9��Ϯ���:���P
�;Q��v��Tp	K��L`��v]���	�,�w�'h��V%fN�i!4�Z캹� V�NLԷN�b�W}9�w���VL���K8!�o8QI����Kp�MM����^�*~q��FW�V�:�/����
��ؚ���RY̟��+y#���;B�Ě%���$�>�:''�G�A��Y�s�cx�j���:'���#��M�P1�|��Q��Y;���m7d�[³�?e��]s�����;+/&���ň�|�u��LL�Ws���}\ȶ��'��"�Sh]]KM2��M��W�Y0��s6U^��҇��ɩ�	���gJර%�ww��<>�STi'H���C��%+�ȓ���}�6;���;hqPD���)�����م`.�J���p}�>�Z@9�'Ck�يa��T�t��x=7w�ř�L�Ee���+B���㯁I���y��jO�P߄<B8��j�R uxΩ �hQWMM�􉋭:&-�U�x�H] ���`@��h
��"�����DP4[����!�t.��R�����a����v�x\�c�:�)�J�(#��0i	��cr��@��#����K+?�XXi��S�%�$��+�ˡ�w"���!��r�װM7ą�;A�CCO�ǁe|<{|�0�Cm2,ġ��2����<!�}Г8"��TD�N4� ś%6��9#!�e�1�c#Iy�u�&<�@N�c^O�&�eg.�$	t��c�cg�^����N�ײ�b��!����0g���$��I �j�oN��5 ���m-���&@��f��	|,G"H���%�1d��$�T��;����j�ݺR�~Yβ��7l_a0g暍��ӕ^`w��
�K�+߄!��;�`��l0S��
�����W���*�}"���Z�7c��͆�HC%\�X4Z� wO�����#�})@Vk'�؊�y�s��������$ʏy���8l�d�K�ζו�˭1���;?V�)r,�>�ԳHX"�d��3*�SwS8��k&W��)��;�����ϫ���p/����)�gMn{�p���BZ�9/�<���8�#:���'��ۭ�!{���.R����5Wۄ��	L����ݾ �� �&�h۳��*Ѹ��+nXD(�f|�	��A��&����$1�?�~b����7f�t�������Y�������Y
O=b�>�h|+)�^��i<Wy�n
�r}L"2S�G��1R]K�YQ��p+(����X����3��'�ʺyWx� %bZ���ŭ(� ާ��P��l	�߈h^��m=2���9t�����P܄m�ɍ$a�~M��T|T!�x `�����3QS�~�%�������4���Id�g����)5Xɖ윹���lT5q�3گ��ѿ�4Q�YSmC�N��~/� ���KcW�r�:���_�����Z�XQ�v_L>ՙFn_D욧'iڕ��K��Wiq�8�,����.���*�8�j�r#�Ӏ���"�`~H�1�~��(T�����E9�fC�MS��U����B��g= �;Q�%�b�E��wh'ޒ�����|�+ñ��C��N�hu��=���)�X�fZ���Y�U�6>C p���$fs3��=���$�@��ɇ����6;D�K\�y�f���d���xq?��/���di��W��یW�&z��t�л!Z3��$�ZXJ��&��j��x���}����mk�
dzy�X%��h�3$?��4�����yu�\��Vq�M�v���M7!��������+��SU�.��+�@e8[�����+��|1�Ga�z��S��u� 'Ȳ�x��T�(l �wm�T�MV;�l7���]�~A")F�����Oh�`z�j+��DN�k���[ħ���U���	E'��`���&�Ϗ�{�Xt_yUY"����360
�F��=�A��;=C�MW�d��$�a?��V��!�SC+Jr+U[O�s^$9yi_'��&�d�^*������.w�\��bB�pJ�7�P!=!�൮��C5�sYSɤ�Fe��pKk�O�tɸU�"x3��[%�0���{="d��ؚ�q����.:�mg�}$.�l�	��^���xi���]�g�j�c�']��4$� �QN\����ˡP��PD�	g�U� o�sf��nS��ӵNUһ��sٜŊ��g k#��\��zpIB/������{���Ây���,ie��<����<0޷#�be��Z��ԕ-"� z�+O���i;������}}�v'��kx�{�e��4;r��O�1N��Q{m�0X,x�8W�\����Ch#m9% ��P}{���^R�K����8ט,K�g1��8@��+�ߤ�	��i�5S���y26�x����af}V+!]y;��M�W�]HL��FRJ����Fn�"���,�U�'��R��Z��Ď�چ�|N{���V��_s�I�ɗ�=�z�<h>�:�	��8��Ԓ�ǥp�G�Q�y��}�����T� (��m���an �v`�3��5,��{Yk[�u�0��-h��
��.�8IQ��w.��gJ�=����p������WC��	�+k��$R�N����XZ��!B��]���w��ð6\Ia~� We��G�6(���(�a/����HK���Ҿ��=@	��W{?CyuG4�0���r�i��y�~N!�E�r�{������U�>�:	n�u�M�H¿i��U:�&�D�h���s��X1�MN7���G��}с���%*�yF�=��YV�K��4����O`���������l�uU]?��.��^�_ ��������~ox��0��P�Hy��Vِ���C��<�@�mP���xx�0����k2�I14��X�Dμ���ʛ��l�/�Dq)tK��Rݖf�����a_�t�o��^'���=7@�ILz�H�e<cy��V&ĵ�@!|�bym�gxdr �}������H_�p1�M��>���B�sbN�6*k�1@�@�7���,\�<0��jK�@�P(�Ķ(��?�-�G�e�j0�l����t ��K.�Ȉ��>}ͿC�}�s9�?�'�=[��(��#9����8O!}�'����� �Cb�⯍�8��g��X��3� �]�-lP���ʺ^�Ⱦ���^/����O�w�@<J��ds�����8�\�cgu&�Ͻ�q%�ȬY�OShʳ)Z�x�d̛�O�a\�'���L��W}M��HNZh�`�Q��N�!�`U���
�9d&`�r�s��PT�vFFp�bûo�hy ��n���q�.Iz���
%���d��G��R8VlG�Խ��1�������H�{�v��O@�J���	�!��Ĳd�}��VR#��>{/U1���%N1�X?��+%;�ўF�Q��wF�e*Dg`*q�{8)�a1�Z��e����5\J�Ըd�: }k"	�IA¨d�������_�,���ί�[���$΋���\V��Խ3��gT�J��m��K�C�x��qo�����7p�i�Q=C+z_�J�,KR��YB�����4��:]�x*��7�ߤ|�H���!�l u������$���L���X0�^����%v %��]�ݳ���q��.Ïg�6Ĭq1�i[FIR~d�i��'�*���������#|O�͛á��������a�Y�M�f�#�Icҋ�x6]Eh�����!8:[z��A�G�mY�lI����.��2�&(":����eܒ�M�)��E0��6�D���e����A���M�ZT��>��:��p_^3O3�V���k�
��h�S.i��:6;�
�����I��g����_!0��^ȥ�^V�-�P8��S���e��H��}�@��	��}��Q��v��o��//G���؛���H'j"�t[Ĩ��-
��|��?C�kNwc,��eӛx�8d�E���u��Z-f�3aZ��}�9��j"$�7� ���̰��׹e�A�~�)��G����i�CS�t��μ�_9̽��c�OG!�;}�h��݁�k^�ֈ�؃X�C�Fӻ ���u�����x
��Z����r�@�����1"�ֿ̜��p� ��x.��&�G�OH�=��;����Kv�Hl����?hM!0-�8s�9��t�F�@�4d�yԠ������刉Zs���~J@�wg8N0s��,Y��o��J���k� r�m���yN(Gn�r�7��2�uTO�Å��<J2o�є�f�����:^�M#?�`�\�F�#��3��طE�o��e�J���կH����27��V��"��>]̋Ӿ5��_��S;U���͸���:k�|�5�"�IV;׷����ij�q-H�ܼ��ˠ�('F �7��JM�����r��L'৻v��7�bj��ʔ�,�Y�Ű���+�<GN�5L,�Q*�<�8��<	��O{�	+�dd��������
�3�{Lq�8 zY[I�NmD�?��yϙ ����� ْz�՝��5��7E� wu���L6�c^ULtHF�F���Jc0b���K uF�X��o��7�y&C�u�N?F˭��,!`D��N����k�DYǩ�����dxA�Z8GndJ�����m/�.��J�Į�����]s9�Rؓ��o<������F�n����9��Fe�7��\�"�Q���TE��V���4�>�4��Z��Ȓs�5�jd'o[�p-��@Ƒ��e_j2 !qb"��C�7Տ�S���=���%��W��&��V�1��N�9`��������5C�(,�����Y<�*c���U��!!�2~�ƴ�O%��A�6�GAa+��R�3md�£FU@A�qRW�4'�" *'�w-�J��K��g���Os�n�M�q�:�P�De�MO����o�g�r�7l�?H�p����+��1����c<ڠ�r���ڽ	� �.��͉���{�+��]+'���ݼ�&}/������<>�����$��L2±@��+<����j��_w�N ՜�i\d���i,�;��ZeM&�� �|#�����]�n��A�p��_n���s4�B�׹��n���(HwG�&�B��&��C,La0���s����\��-d�3�*?n��;�C�j#��A���&.p4�mQ��2��؂S��SyE�L��Hn�G�F��o���{H�]4�	��Z��F��X��˛	�t����EVF=��*o���F��o�n�$w̰�焕�e)�R����ϊ��l�"�����X$�M��ه��� �V��u<g2��9va7V���<=�9�{=Jŗ;$d/�@�:7瘺��SR�1��C��GY�=�֮j\>�L�V�^���C���b��z�ة���+/p�.�A�<��lFF��}qN{��pfR��x}wwq�L�������#�ΣO9��˫��1�@܍W��ܦ�,�O�cU]��NEk�r�L���(v�)� $�������pLH�v\[5{/�GQ���.K����VC�e���.����,�� ���f�\�$~�	�gɴ�8���-2:��N̳l���r!��\�~NZ�µP����RL+Z��~c�l�/	���*���V��*G���|�8��ޏas`��E/Y�cWVț!��gD��'MF�>D��Z&��y*e@,X�xGN�9d�6���3��f)�;�e� �J���ҕq��ML���%���K�V�H�~�BF�����D��ܑL'Zq_�}v%�s�H�:ǆ����'��^fI�x�a]6��;�"�������%��N�7)�"�mo�t�X2��Oڵ>�$)Y#�ky*��=w���0�9ʤ�E�lK�����L*��[�K�S�5�R[CM{�;aAK�d�qf\��k�ԼLz��Uy=��;�웽�I�6���Een�D�J!�ߘ�x�M&��>���)�S�������Fj���������IgQ�V/���oe�^���M`jɕ�r���UIM��6̈����W����u�:�E�;���[�Pd<bdQ�}G(3�8��s��`*"��B�JՃ��ȱ4}ΟXE�4�ĴŪ�� �W��u��2�E����?��D�]e-��b��gLF��T�����&�#Grb�K��-뼔����U�T5@����m���"��g�=����[�pDz��y��U7��b펷�����D�\�J�������yFi�!��Voy鐦�>��5�I�UK`�T���I�#?C��W����@&A���8t������S�� H��N�˲�����3������3�i����Awa5:x�v�HLŃ
*�B9��dge�*c��]�UG�%U����Daw�)�7�j%8�G�!(��LYq�����?R���Ss�������]h�L7�%टR���OU��m�(��`qc�A�ml�	G*2��4k̒#
��<To��l{K��3	$_�dCU�i"o��:����n��&-3����#�$!$��!��˂G�I��~x�s�.�m˃J"��P�yD������R�>���D,⹡��G'��|%݃^�A�T$�X��D�0}����e=����GЬ�Ijh$05>G�LxH$��S��Tg}�Y����@?�������ކ�$!�I�Y̌��3I�
̓�:0�H�~�|�Jg<��i�=Ees�8��RFFbB��a�O����+Q���SB�����fK EB*�lL2*��ŕ�⫩������yr�c�e9f�i��jh������4�2���xm�G� �H�i��臉�+��وc�9���9�����[�����f����tw;���co�q��#�R�b�Y�zOv����T���fA�~��!��t�!b��c�N��`E�	"j{��V�#�}i��".!j�����ʡA	F��8Xz�	?G�5�L��'��i���/#�9ǿ��q7�VU3x���˼35�i�|���tE��+�h��vk������`\F�Ǔu�]rC��X���`/1�¯�dˆ��mA���EX�=�Σn���&~���{/��[j�WRn��_4�4���0;h	Ma�`6���eϟ臺*M��k��6�l�q6�����廢��qs*�MМ��S'�%��7Q]�����	����7���XέiD�D�mQ]L��k�ê�8s�����έ�C/�ce��HUv,~�g,���ڮxz�bk3�ʠ%�,,��V��<�ܒ ��w[4�~9��;��Ի�	-���b5gx�m���L��^�5���AZ Iּ٤�&,���X�r�Y���uPy��hU/�y�٧R�F����nF���H�q8��#e?︶��AUZ]V�eUD�� lxyͱ5�������P-��WN�P��qӞ��.d��P���������H��S�G/�Y�e�����>�(r��i�W�_,�x�iLS�ϓn��B��?�s�cnA������S�
�m�����U3O�l�\P�I����<�ƥ�oU�Wr���֊E0��ƾ�	]O�d�G).��A�"
�K#���L�7J�j;ȣ}��ْt%�����^��|"U8U�.l�^���;�O~
�=�^��&��w��/O*�:��B|b��V�d-�y0y�Ab���k�,�sBo-=G�&a�����s�_� ��.j٪���L�*p���Z�#�}�ky R���$fF���*�Ɲ	����t�{Ηga1�Ӫ�c��+��4�1g������XO,&��3o5TPIo�d>x*��$QG5��f<����\�IO��	�)@,��L�,��X�BE#��*U����A�>B��{���!�y�λ��Q�6$�6w�_,Gn�Sd�"�������Am��zH���14�iD�E��3�v��Yd���NN�Zf���z
P���b���e ��1eQ��Cnq	Y��1��$�R�ɪ�0���*z��V}�oS"���+�}�n��h8�N���?���(9ԧ�x���~�:���|�ܳ����'�ñ+H�����'���^�����$R�5W=r5����<�r_�4��/�K���#�E7�墴pU�J�����`�ړT`�I�� @۵\�u�ţ�Gb^G8�n��>X�b��mU7����QU& 6~0m��fr\7À,�0΢�t��ʧ�x���(0�8�ˏ����O)Z�a^*�5S��zxv�Vb>[W˷�+�K��eѐØ_�^�!�@m<]�Cc�"�*���=�e*�"�F��?��I`�ь�L���͉��)9Z���GLvޒ�H����~W-��5�pI`c��Y�$-b�b˓Żܭ�=��C�{�fus�@�{�nP  P�p�����oeI~�ܡ���B�'z����5�JR��V5�B'��}�|���O��z�4���"��� v�;��i�Kr-<���G���7��Ll�-~�(�38��feO1����p8nd��^��΅r�Ѐ���X�<iW��6h�Ϝ<|$�D4"?h�mꪫ�2Y�=�d�&��&�A��¬.~+��|���%i$sQ�9�r��e�J����Pd���C�����Θ>�����& ���� ��/���s�i�V�v�N-��TG7���G���ɮ"�J!���֊��e�K��Q��è�8^~ �J:b�f��Td�)f����7e�&E(zW��5�2�k������,��`�	�J'~�kJ�:o	\bH���2[=Ga���B^�iLz�kZ����B[�����p�)'ej�OZ���HpCs��!�ư#�Y'�[���򡻜U�aI�G'�����ܺ���Qx�s9�$C����C��0�2���� �f���-�wd�h6��9!�����m��25�w��]�)l���j��ɨ���dõۗ$�7foF�,;��$�\�<�}�3���w#N�9V��c����,^�[|Q�C�GU~+L=n�T³� \��k��0��z�����D2*�����A�c�*1��d)��.QҪ��:��|��5��w�dm�Z�+�⋅����7uB*|5$�f�9ћOz�&Q�߭�jx#@��d/ݹ|��B��!�s��f��{�E�ev��>3����d Њ�z�A��E��lu��3aS(��쯉�m?��H�]#���w.&!�#��%��B��!xU`;&O87	�o?喽�)��e�7`�?Z(�k�`�f�_�����څt�1ll��}�eT~�f���jB7�ns��E"��|����hN�N��$pe!�D�8�U�\��#�}���b�g;�Or,�r
��Ǡ�i�yH�]ZY�1]�S�*���{ɡ.�. �W�Elkc ؑ� k*���e4C�K��p����]�/�������r\�ɧ�K��5��:j��>e�Ł��ܩv��S�_�'��,ƙCx_���EIy�ڽ�hm�����/��uZ���%P�n1�u��2� ��`��r2��]B̺e}�0�y��'��W0گc������$*���2rN�_�Q=c�<��pϯ�ˣG��t���"�Q:�7#�Ͽ��
I��%aFc�0�iwN[�J��Q?B�+	9�p��7���"� �6d�*�QQ��n=�v��@N;����no�t�ϧ|��`�������Kp����d�+�����s��F��5q�c�K?�E(|��ј�
O/#t�A��֖�h�L9)�Q�63P�����Zn��yӾ�<,_���.���p3�D��[!�H:׶oJ���5��t��bȄ����9d}�a[֐ئ�U�5x��u7����ݫ���ΎRe$4l��C3P�^K��.����N,�7��C˱*He�<�اj���pBE�F�%���[\j+ ��2�l����j���~n~ɇRH�y���4~�o|���o�N2���l�,dQ1������D��2���4��hd�zف�T"�v"���{ϡ��;m_N/�|L`J�f���IL@�tw�+���x0�k���2�6�����v����71�t`;�˒�@���,��kU��'�#�#��c�L�;���H���E�����?C*���u:��:x�����ܯ+W���ۘ�R3Q7O�_r��k���o�!��^�}���Ρ)��YJrS�SX�ts��6q�ѹUMLY��u%��l;`O_�+'�r
q��0	���u �q�;�O-����M�8�Qwğ�:���Rv��S�dh	ux�������g:9\�A�������1]�@�Y`�_g��t�)�X��u[ 5k5x���ؤ^�����@M�������>U��w��2Ɯo��f��&�'��/�@H""ڕ2T���� L��p!0{��8�g����4"b٭R�k��pN}z��x��J����]�]��M��*�a0�{M�.������!�%/(<�η��4���Z�?���([��KO��}�B	�_�F�>�d����ȋ�K��:w�;�u3�7����rꅧϦ@�ab{��u��UN�P�u������ॠ�t �n��I���\��L�#\.凫�%����L�L<��G2s���]u��ϸ���g�G�Q�	�N� ��Gb
r� ���0��Ůhć9�	�A�Q�Ƽ���Z㵊9L���k@��mHs"�|Yu�����d�_~���u�m!x>����� ��M׎��N�P}<ED�0�����:y�n���S�F;��.�^��r�?,%�{d�Ll�ܑ7E��XB�8s�+�Ӣ�j�g�W>@�y��8D�>t��������ެ���G^MM�o�K.��G2�[Po��:���z6{�rs�/�k�\�^��������q8�욣�@�s� _?�B��\j!�Q&}��bC�����"���9�MꞭ�KHX��"wl=23)��kg��_�J�‾~?� P�L�Ih1����9�j|���c���+�ˉ����ӱfF����fm	z��Ut�,	t|���)S`���7¤)lQ�m���̈]*Ё)��t���y�&7���_SC�1凤ʧ �+�ڭd�Y>A��Q�y���D����b��n��������cM�Ħ���o��m���Cs@d��_����jĥnԓ�JF9\:���?׾�Z�$|����������1�'A��0"�4���񓿄��wXc;��<�~3w�����u�~�AΒ���}P�֡z�l)y�ހ�rZ0�VFb����k�8�N���ǳ�K���Lxڣgj��6�1� U���4+�XWl"�D&���5~�'c�aNw
vQ�h��=�ìۜT%D��A��3�S���%�[)^� �4X��V �<�XE�3�s��*��v=�7}e�B��q�շD����By�H�����4�����v�X7d���6G�)��r#�c�;�6O�5oJ6������ɝ4�|?48�/!�Ȭ�)� ������K�jߝ˟f���}�&A/3��B�u_(�'ak��_r[H�9���߱���u�x���ҭ�<������c*�#��$a-؈���4���N�6{K�1���A����Ҁ�}��Mg�R�8�)a�U�F�J°�������*B���V�2/A�=�1�ˡ60�%��a�������䓙���(��3܎���<��!0i\��Ն��J��,##�`�"��j��U�=OG�,I��C�ι9/������yw�"��f����2�,.���^2�Ju�E ����BTQH��rb��`�F}�lC�l��;f�z�VQ��/_�hu.��_��B���-rl������jot�L�ހ:���ȁ��fE���{��g1&еL�}+x�\�(�( ��ť\fE��Hܵ���[��6ə��#�6S")>�5��%�@SꓔM��l:o��@�����+x�mpo��URBDL_��|�ƿJ,2b��Y�M X����;n�R
���c����)�k����QR�8�,�������/���4�(�{��:�����n+�8:�o����Ǩ�`֫�X��z�)xguY���=���,h��@�{`IX*v��]R������?��'H5�>n���� |BQiw����M���a��$m�J��s���J�v���2Ý���*�סE+���@�*-|\X��})-[F	�PIX �f_~������:TզU'I�,��:l�ƚ/8�	~�{;�`�M^X��,��(Zŉ #����/�j�hx��b`�+�Y▓��>�E�-�����l>'��p��?��k�X�[��4�j���>|����ޅd?��8���lc٧�)5R+/�Cԫ�����!]�"S:&Ϥ9X�S�h��'7b��BC��`*����8CJ)��%V2���9����t��� �q�\'�<��5���6��x�{�9�X�������$S�mU=���E��_������?�&E�C���x�7R6�Y���D��ST�w�j�g������5h=,�Ǎ��
=��>h��?6c��v�`����,�_�ibX����]��+
lu��4j���˥������+�y:pJ������~�|;�sn����N��N�%V��{c@�2����!� ��Y�=�����0"��k�/��y�J�
S�I�	��qu���fq��h�l�5��@W�L\�*��#�Y��H�ث�kR>�ۨ����U6�lc.ޕ�����m���CT	�m�-�x�Ԡ-��!����:��7gTۀ�����~ݭw�Y~ԩ�j�\zBA|i�!_��4��I%���/;N`l�9ײ��I�\��S�e���5���)M�3�7�||k��ǻ��fU���z�'�(�4_.)~�Y
�@g'��t����ܤTo��?G�`C���&o�&�c9�sqWP�D���^o��b,�.��w��>jMl����o���6,B������l(,�^���H�����:�xVt�Y�e�ޕ�&i�I2!�6��s�����n�q��T��1���T[i�rE	���. ��6e�a������t]k�ΌX����9��1z���@�CzϹ����u��Α?]s�0��"y8gNC�d�����~��b�������N� ���ؚ���/�Q��>tA��s4���c�e��U|���b�>&S����å�`�QO:@C)Y���0q`��֌pNW�ʴE�v��+���A�7 �fA<���5�1�!�I#'^�'�1v{%�-e�����_\�^�l�����d�	��>��j�0;�v�w�:\�_J�㑙B����E��,>ذ^w؀��o�j��rsޅ.
�E�}b�r<�����_���9�4=Eǜ���X�o3?�/�	�87z���8X����#� �Vl{�z\D�ԝ�M�R���R��C���� �jO��{��#����=7l]Qj(�]��n��hp{S�
u�W��
�+��QW?���3Ӌ�ذd��UX�β��%5�x�dS�ڋ�#E����T�����f�F�Sa{�l��v���@�y�n�m,�|7|�	#�:O7!f�@��{h�s�&����A�k��^>L@��_�^����Do��f;F�)s?�#�'P���R�ꯛd<R]�D=�G��n��z�2\p�+����㏶�aPH~�A3�F���,��q����4CR㒆y�)�HeM��Y��G8J��5�D�x���R]�\f�0��R��ہrc�����F���X7�໿���5��3D�hp,"L?,<��cR��BUv~˩vl(7J�7i�W��V,�7'�߲��W�����^89�(l�D2� T�4�E[g^�B��#���f�H��P�C��s_�	��f��ң��z����8V���P�S����צF�H.X�� y���S�<�UX;"Q��>�_R�����y��,`�&DI1A#m>���䂧mԼ����̛E)�o��ߩP�)��ݠ ��R�'w�Q{�u�*m�3
�4��
\�E���"��ğ�%ͭ���@d6�6a���
�s��d���Zl�@oO@�%t���K=Ujd��ƉN�6�sD䷒�q �å��~�"�'� ��e����KK0O�_"�>�[!���o��-��.��T��e#x^(��-����Գc�{dUw���=ɶ�dh��h[[�~Y���j������Ј���?�)��37��=�gG7���1.��|��P+c�qo*�)M,�5��E<2Sg����}�}Kn�gW�z!����\��HK:�q�Kn@�F(G
�c�-�����IV�=������N��C�y`�>z�V�׃��kD伛P'Z��}�F���Rr��==�O���H�W``R�L��O�̄�O۬��"��CfyFa�Ƞa-�ޜ5�Jg�H��p��D~XC�g��:� �aYE�q�^�ѓ��i N�e�������y�*)��ԅ�h���W<9�fH�%�cG�JS����;�R,+ܶ�7��Bu釔a}�(Mg���3��ڇy;L��&���+�kź��K Y����g�;qK�<���|3��g�C昫Ӂ�Mv�"*�׳�0^�M�|��C��!��H1��e,ۇ�p���ɯ�	~s��k�f%fM��b4�s�8�Vp!97Nk1��_�p|E���M�:��_�<��G��d~p8B���
Xo���M^��j�k/'u�c��1�W7-@�!�X�$Q���yD�u�I\(���DMl�����\0�B�k���N�O�Dm�3�~n��� ��gnqϓ�|V��k��]�sظr�Z��ѹ%�J�6��#P��g�i�k��(탳����`]�ݛ��LU��w"b�FE�vg��:f�w����Ԯ�k�Dtƭ���-�O�8`y���(��U$\n�8U��O	F��p&i�0�7��MP�j	(%����_)ml�<J��v�I �Qz�(GPR�Ϻ&u� ۀ�`�cX�]���+�j�N����@�J}�j;���u�����Z+k������Z"��'G_QˤҾ�����s'�-Դi����|�?��Fώ���|�����N+��}d3��$"�}/�o��=G�\� s�$�*n�e3�}��ӕ�g��hu'}�j��em��5'�Z���y�M��I��?�5�M BC����9p���T�E�<�����m���=�f������A�i .*ʏ��+d�u��jE�'������9P	�#^4@N�:�u��.�a�F�8U����Y=:	����&O�%Q"'bю��[���9��.��R �Dɳp� �ܠ�7��G���^ ��TT��>���'�0�X�N
�����Ae55���thف͑��f_�{)߾	�2(�ˌ����w.��z!�PX�MF����i|6A�M1z;c�\�ћ��1�?�����X��g����K���X��Jf�|���B�&~tPm{�P���@]>1W�l@j�D%��g  A6�����\(|��B�W)�~ j/K"#�s�ڏ˳�	_3��0�]WV6&Т66�G2z�aP���4\�*��PS� �p�rsQt�
!d)��0�8�H��%��c�*�?�,���l�b�%%�/y�?�Tpjr�K�/G��	��t)C���K`�%�1{��_��~8��q���M��O����o�Q���玳>�-Ef�=Ƈ�������c�>Z�|+�l4��7�+�|�ڈ��=+f���J�spOಸ���)�3�V��v�\��7��v�QW�J���0��[�5��TO�����\RkK�#Kխ��r��pQ�W�ϖ�*����?�e̫�tt=���}�]���	��zl$�&(�b�bp[�3\��܌'��>�Q���M�ʒ��,�H3� a�G��e�����⣉z�.�y+;��"�#H�2w�)iw#�-�$�opߴ�8<��]*�/g�
�Ӟ�k�+�}9�_~��U�%u~��#�Vc���'����?��!���k6�F�MM����f�������ׄxY�{$��ž�C)��vM^�"�JLy#1��7l���3"Z&�њ�,Tp&Hg�3F{�n|�E$�u�t �E��T�ѐ:��"��M��!��R���|ׁ�?ϸ���ػҌD����{n��z_��9�v��%�X�7$�K�ޗ�3R'�4uv����r�+��9k��zZ��ϱ6��$� Y�b��{\�7��|�����o�ݼQ�����E��2)ᾷ��N�ի�v�az
B)�B�o=-��1՚Hm�m��)�`�ƸH�.G֗���\Z�MO��B����	����eέ9ھ�(5[}�Jݦ�D��ʻ�E��B��jIhI1m���{�CRo8�"&�g�Ļ���*aE7G��%p[wa5ݾt�
y���ߔ\:����0� �%J���3��ۡ�����N@�g~�>ڬ��o[|wzܲ`k�9��k~����2���*�ӌߜ�G)bv���m7ɾ�٤��nH�0�~w���]�o�@���<0�$�ș���&x�����(c�H�Q�`�;d���� +�*�@	#�r,�Sg���.=u?W7����
͈���H� ����N_��;������Ҳ�(q�'�NӺ��࡙
ݱeE���������-�?����m^�����d��k���a��^���.ȱ9\,?<�s3�z���_�~L^t^�py��- ���E�E���b!Ξ���I9��PMmw�)
�4��xu�n�WPզ/��+��K�{��WC�B����C��#�:�$�+��~��=v	�H?�E=:¤�p|�&��#�kDF��A��OC�W�8¸��~x��5��J��=��ʒ<�6}�{(ҩ�z�ej�`�R�_+h��Q��~�&	3P2�>�^�g��5[�����Eo��B�Yt���Y�I�|�/JH{�_�RN���0�����6���]T��!�E]J!O��g�lm��C�g�I���<O7�l�fBOM����`Y�X�8�5�~����*��aMc�D�tc�L�I���S��g��<�����UTP-Mj��kN�~��/j&�ö��R�V`���T7�,5�!)���"����ö�xDK6�T��kt�(�_�f6p������x�G��N/�$璎Hp��	~o����|~5~��(4�}{<by֗`v��>��&_<��Vq��,�Z���B�uFS�|Bx&��8��E?>��4!1�居꙳�����ܚ�f�fr�9?S���V��-ӈ%��b��&�lL<�(b�ox/��#"�I�{��[tg|,LIO�p��j�Gp�7!�h��� ���ʥ��[����`�aH^�kg��89 H���̉�W�»|�Il�ܹ��'fs�D �ɍ*�Fb��"Y��µ?��f�v��	#�7�'q��4�_�[�η[j#B׳߿3�R(��|]�����i�Vo�Q4��N5����z2���PFQ��Ȓ�(���Fq���U����4H�$���$���[���.��g�4H�����a�����a�g��IsQ�H#q��0WnIiY�q�ݽ���r�!����&�O��Q�L+v���{N��AP�2$�j�{v8%~����?�ͱ���)P��u���iS�Z�`���1�,I��2�>�c����M�^�	�<7��+qrf:�D!�ɤ����n�x&wO���)�6�l���L�����6�Ӕ�ͪ�-�����-�I|��&j��0q�fI��F{�y������*�vf�r��E���_1a$��� Yr(s ~��G�Amj
�́�@w8�7�
�	�y�l��^ep��=�~I�"�[��\�0Z�x�>:���Ac��TwY�L�B��'N�-.'���GF��M@*y84NE^��1���	��k������J�^��:��3�C��B��k���me�A�Sb%X�fU����}�˗�� ��1�o� 'u�xY��6�;��f7ۑ��i��
0ا1g0�~��6�ǟ�����(���kP�o3O�1<�s���c�Ы&�JNN4%^,,ΪsO�r�2u� �{�t�tE*;��@wMD�9��E
a7���c�(O���������p,��^1��L?�<9u��[ի
@�."��G	V��,~r��A1bW���$�{I�ao��w	���h�(C��}#X��2(�Y_$ݗ˭�w@�e��K�?M����\�?��zU������Wk؃{�cǭU]����5�����5���}�3�����?/g
x��P��̹ ��vo5*��7D1���N^A���B�!�ٿ_�W�ӛ��p�Ԙi���<�j�X��;	�t�x��;�z���B+:iN�8u���=��A@�������m>Z�׵�+�x��o00Qs�^�YR��"��Dr<�u��g�L�9�h)�^�F8d�?��_�|&���S�1^C�:�T[~]��P�+&	�W��Ŵ�aPנ������,��&Z@�Ǘ��"2|aJ�)$B#�|�2q|����P�$���$�e`��#��w�{�iY�p�,�ƹ��5��3na�NP����y����ơ�K�r]��0-�}���_��o9�����h��ѕ���$7ϖ���w07�H�*嗁�%�[�T?�16���װ��N`���NvdC�'��
w�2��ՑL��6[����weA�e��/:@}���*��ĔS�5���:6`.wGwz9+���c��W�~Qn�?�<����'�.*]�Л�$x�4�uW��w���:�0c�:�����_���@��hB��V;���Iڍ�Ԏ3�
�}�Xh`�ۻ�_=�Q�?i��щQ]�)����ߏ�>,]�'��w(5��w}�Py7y��=��~x��%�I`��_�R�
Wk(����B"���<usL�So4~g6�q�=���4��謘������z��@�N��ϯ�)�-�)n���8���/�1�{W7M��b�f�4���Ö�p��D��}�	��@F´�=��v���q޽zs J��T����="�A<J
u���QM�1�2û���!�/*'�Dk~\Y�2'��[w���Q��p1а�S����J�l���~^����ty*��Nd���E} ��O�:�ZFlq܇NV��Hl(���-���}�:�p5՟�ʒ.]�[�s�h ���Ca(P`?ڦ�)l��h�h%9H�����x��kcƬ��Ljܝ�I�s����+M���ۚ��� S.r�t�&|��7, � �́Sw�i�!��<G��3�RK�]u�+Gf���KS�ue=r��?��)Q("�^�ժ�q���c��:��rn�M*uv6��q�4�c<�"�ѓ)��'���#{�����!
)j�`�0�-�Y�S,�iF��jW�z��~g�_�P=�]��̤J�RZ��,Bge�)��A�٧c�5/���Qj��=�i1���� ��.�?.Dn;�9VO ב�R%�i|��5`������ -�?�K���1�,dy�i3�OX!!�7��5���B�;:f��س�^�'�;�տ��qLtY�ɹ��&"S�5_��/��\��Ol��ZH�(��S�"���/��LX��K`�G���6�[߬�ͬ�P5_���z�I[�ͦHLi~n�6i;�Imz�l<j!�,
c��YH���a�E��f^Q�)��ϐQ2���w�,K7�].��$ȤR��S)c_�y�;���-HD{�g<  ����^Tǆ�ޝ�r����N*pH�ɮ���SCw�娌_�8�X=���ID��'�~�fYG\[:��>f��s��qM킽��ss��ch�湞ucP��.�<l�L��$�v4l�|��h 㢉�Ӊa
�%�"��4U1��%8�N=�ne��]lczR�ݠ�����3��Z��)W=� /�"�I,=e"Wz\�(8dF�|�d&�pt�@�d��o���>�|��I��a̾`��{�'ݤ�p��a�����te>ƟVz;��u�5S�@��LZxB6���T� m���^�R�=�Ê���"#�6��dU1����fh���d�:z���!_��)wNj�J!�S�x���J�KXagE2)�0��ט�ъ�UدM@�)ZmM���[�˶t����s�*pq���{�wXv��ϴ��$�������E��mū��6�4�A}��j��AH�D��J�8S��V8�[����L��q1B6K���X%d�L-t�%�K/�^�f�p���?b�Nyx|r�/�|x*SX�C��.AH��\O_��v�#Z��ʲ������S ��G���%�1U��d��/���>2�}��<�o0�T��ףzu%C�4��[�k����p���љ�/#�eenE|�W	)��%U��iA��TLO@��'�_J�H$�v1��Z�0��|B�~����)
��2麓�g}�1[D.z��_����k_R7�u�ٳ�l-�{H�F��s����-�#=�1ƆР��ï�3�I�,z �8J����ǄkB!kk8���dl}0�����>�=��jB�d#�_<�e2�4��?Z��4�(k��=?�w}s�e7.%x��d���?���Kt�_���L��_�-�ZH�:+-��\�K�-�`�	[�F94�<"�8��"qcn�߭�ȧ��7v}�)׉R�;��j��b[%��d�R�Ox�x1��O�<��	\�0�Ϻ�w� �!=�Z���fy�3ȩ�	�aX-�6��3�7�~+c�0�����]����fA����~9?g�?|�]�\,
?m���إLڤ!�i�Au�L��#
���?�|X��Bzf?p�}g�3w�ER�`T��f@�RB�:ʾNf%���%��iY�*��� ��t��K-�T�d�l	��_l*R�D�B`1'l[sE���a-��g�/غ:Ho�lo��V) �k�_	��7�c�7�yЛ��w2�ɧ�У�R�iRs �@O��u�j]a2T�/@ F@5����Ґ���u��.��4if�Y����Ajmj��20�bH��r���?���`�߬'`&��a���Q\�������paǟi���_�pɡ������e+"�ܲw7�ԗțS2rm+\`�-��eN��d)Y5��5Cז���4O�w%��fz4%!�r���O�K��FS�JM�ovջ�%��;�.B.��5Q��n"+��l��"�j±I��n�*��p����#a�Z�)Kb=���'�0S.G�C]<0`���	�p^��S�z��7\�Hz�VI����Jt��j�	��"�d��;H}��Z�s�|9��kK0�c����Y	�&�v؏ʦ�e���|b�o;>gego�UT��l��?��c��L��K����O�
��t�{�5�8�89Du	���A@����V{<��5���ǷB,�\�(mU[~m��E�W��o~
ٝY�X��I���;���5�Ng����{��zuR?��s�`����c~��3��d&>�I�'�5>�>��?o��:����͡��C�"ѧ.ć�Lgk��>�T��ݤ�uUr]ħc�*��� !G�"GB��M��&{(� ��,B�
��HZXT ��2!���&g��"S����)#hO�
j���}&��R�8�,#'��素���CȽɬ&����v��B�G���*a1����g{��	�0���HBF�ޜ$�j�7we����I�ҳԱj�!]�8���I�.� =߈\|�9N}�>g=��~"6ǯ9]zk3E�:Dsh�/��J.؏0�k����	v�/��)�8��8g~�k�,kDh\C�p���$��B��W��{}��G}�p�����裃�4��O���>J�$����h=�Pʗ�T"��{��e��w�|�;�K�M?o��yT�d�1����\8ņ�f�sL���α7m��0��3w���k/��*E�|����,/����.��i-\�`��z.�$%hV?��]HZ��	E��?X�8���9�j蜯�D�KI��ȮM�#��L4>�"�H��%�K�όSۈu�i�j��8���6�i\���N@��@�zBo^Iv�CO�w��=>�C�i_$ӟ���S<X�t��TpT�o^x��2�e�y�W�3��T�}��?�~{���S�β|�2 ܇�1�����>x#���E���%�:���8Dh�J���k ���9���ً�J"^��> Il���k �N�����4�a�4��,�F"�8����0���ӳ�T��o6���yv��^�D�u@s�x��'�ܮ���Fq��T�,J?�I����~�h]V&`��'7���!�V��Wb5�ʂ3)H]�:H`X��M�i�FumFs��8��+m���%?f��	��H����[�$�.+�-쬼�Ln�EUa�8m��8���y�P�l%:�65W#�TW� !���`SS��d�xr�Ň�#|�����H���!II�Ah�Q�k�����펆U�i�(NiU��ך��f�9����Z�<�<|�5VU�h��ʕ��\I��A9Ԋ�<C�
9@�g��39)?���f��w_��#n*h6�4w{7K��d�8r��l�Y���ml�6��Cäkp��I����#I�吤�z5P��6���/-�L`z߁$�T�T����K��t�b�0�<)9Ƥ���ǞKw��e�Y�*2�L�nħu*���j�lI��s4��c~sr(�6��,v����ӂF��������i��B�}}��c�M�逸H�K__���B��GV��Yg�Ġ4�`�MS��'W}�>�����N.y�,��vZ��0����q�����,ɇO���0�]ɰ6��ޮIw<�c1�F�kR{|�q��%���T���^S0F�|t��h�������嬗���\�}@K��<�l�%�3U-X�k�x��|!r�܂^�f�\�|�9>�B�k�O"���lX�s8�0��)�#G�P�d��~T�b;x�o�j� �]���m�:��·7�Hm�d�j@T_r�b�U+%�װ�pv������E�P�eR��ƒ��0�x 	�ÈK�y�Ui;?I�;�����&�@۳M��-�[���� ��9��(NŚ���f���Ŗ����p�\r���=s��&�:@�oZ*�/��~�|��[�/U��6�d$E�'iPt?�J����v�	�j媊��O(0�lHP��4�Z�g�z��!J��rG6�F��R�5��<J�	V���ѲK@�s{&�?� o���iw�p#XU5� |�Vٴ��O7���[�F�����ۢZd9��;�E��~}��ښ����=r:�œ4p� r�Ė��G-U�IZ�.4H��s�!��>�c�*�pդY����]�rnǅ�����7VV�u�U��'1+32lB���1"r�&%�MK��mP������K�v��~��#���N�L�X�.+��h]��Ὅ@���[�'�f�3�W5�������``D��_��E��]��.g��Tp A��%�tm�s~w:څ�1�b���\�S����&�������֬�c�Qp���fmo#���i�^���(�؈z
�"�6.�Re�!�2���5�`f&t��^��~�\�����.3�$�I9!�HM��݀	��VX�RG�C�I����P��C�3<�۝�Zjo�VLf��+Qݳ:`�f�X�Y��%G��ߠ6�)��
��f��KF�0������R���wsR��n��P�3�q"Jq2R����(Q��ce����gR����UZ=P�0�4 ����M�	&f��l����u�"
�4�8�)W�-����;I���I}	F1[i^8���<	��~��|U��Z��y	��Vv?�$\���	���X�gk	���
�6�o�]$ה�d�w�%��>q��ڥ>�=*	���A"�̙	�dǙg�S��eh���ڔ\�]���.o��_�D#�M.�7�ҙ�Yv ��3tB��ݤf0�q!�����s�{Φk'���Z�A���5;���m�`���
;R���T7/�H�ir�e��_�O-�*���d+)k���Rf�G��ڨH����J�Y̐�G�����ܑ�<\��i���T%q5X!	������TS�[����	0_�v��(�:M��ȸ���59W���S��l��Dĥ�xK-P�"��+l�y�  �o�@ZI�[&�kxȔ��ٮ���4���"[MPtC��[�X��y+�"C�S��n�"~��?����½���^Y?�>�c�r������g�k� oFhD3�TK��"Z��*�c�FG�f�V��Q�h�P�����A��?x�d�T�&t�R�αaм��|�8O�� |�B�<y�T��ov�O,p�~�SJN~�Ő�@òs+oj���+"HU@�f�Sg>;N�ڠ՜q�F�4�����T�3)�]��Ơv=b���c�2�N�E�\��:6�<�fv��������%��Ƿø�`⮒��h��{H<�ōb6޵n WK��N��H��l��0ǭ�n�wUϡT���r�_�Q��Q�K�ee��.��}|l��yS�Ы�o ;�R�oɧ�k��X�4�?ۮ�\	���U_=�3�FH�sϳ��s軌����>�5W�猳��w����:����z�)�*���%)��z���%o�}���6�e��B��
�b�U)Z�*텛��s����A�� b��ey�tܦ���mSp�H��%7���M�74�]U�R����h�)�qU�[d�Y��w5)��m�`���+[GY�p��n�9����ܢ�x�Jj��K,t�X8��]�&�;�E���zao��![�%a�D.�Wm��1�r�{	�ʭz�O.���ȹ^߯VZ�J�D���צ`�*�e��9�.?\�_	���Z����}����w]�f��5��(CRX��@�{����`�N_���(g�)p.��s.	޶���e���pO �>W�x|R�2���*�W(6ϰٰ]Ɔ���@����x�cSy3s��� FT���gyL�!%���I�;�τ�	�K�G��M���iI�''�_��:&�Y�nW�������o���nX\,���yj�v]d@7U����W���,"�aB��W� 0���X�Dwv^L��F7���kr'��K�����l�8�ǸXY���o�ذd��$�9@�I��$(�C��bc��/�9���u�?#��yi����E��= H����A�?�'�{�G����9��S[�2��֮����[��LVti8�Fh[ң4�3j��z2�/v�q�遌�4�p"V��<�� �iNHX�a�hr�'>����l|eY�?b긜yCJͫ��/h��t�5P�M��?����5胫c��ǜj�����ln:��u%���ӂ�:b���鿮a��!���A!��z��«�z@���f$��I%>(oVx����c���z�����j"@�H�����g����7׺[mE1m�|07>��@hoh�K���+�,�6�d�s�An94�N�)�xY�ʎ3)9�ڪ���w͏�I]9qx�<�n�7��e�3.��.=OTe��fd�騰UC�������<�}`񂪂��D&�UQU��Èj#�I4���F�F����Z�7s��:N� ��K���kQ+^f�B-���9�Dl�Zd&���cN)�hL!F\����/�p����\��F4#�V�vHoB[5A�y�2�$l���	��1~ ��)ӂ�Q=�[�Hȵ��؆��)/fk�	3�\���.���d%o؀�a��'�=���F���-%��u/�>�3;5	�N�G��(��Wxi� �>mMh\�7�V����?\> W��>,���T�Z�F����R�/���K�l�{�qj���\��T���Z��];��|�)1��Z�F�~�JQT<>:��(1�-i����auw�d����wmf�w_�)�	T��\�ޑ�o,R.�n���l�����X|ߓk�^��BH-�r�o������df���C�mD��fE��5A�a򱷌�]��ױ>(�CW�<e�huR[^5"�qu�Ih��%��;t����� ���'d�������6�/�?��`�X����g.B�'.i�R�d�k����Y֪4�p����}�oio��� \��@<��Z��a��#��x�:Q�Pfÿ��S�R,���o�Qh<�S�?�� �ؖ�@�S�eVL>Q���=�wy~	���1��Ӑs�(�<=
H
<��`�V&��Gp'_��A����)c�&�1ܾ�D�&��&�}4Z��wKڼ�Z�UN-��2|�*�P?+6����
���VM�[�P���BơG>Э���\����2�؉	�NV��9rh�ȧ�p�BG/:���H�����}�d�W%ڒ�����!��f���{�¹X���J�q���c5�E��#+#<6�u��wI����Ex�Ord��=��/H4J�N�ݦ`S��"��� ����8�l�y��F&�9m���ވBx���AqOU���tl�Wͳ	�>��A�����t��[�6�ʏt8�R�ޟjG�61Ρ�w��l�+W���G{aN�*�[	ۜ�K�P6��*MR�X.�-AW��c@D�jJJ�ϝ�ĔM�<�L��\������P���-+Ky�o���p�hi-�T��'��,����㙫��n�*����E��3�+����/���h�?��]�kVy(�ŋ5�-��]lT���R�<.���閴 YA�D�ƇsgX��P܉�������]r|�z�a� trp};�O�����І@�f��I�"�q4oJ�6
�+��9H8�:g��Fv�)����?f��k����%�&e)���I�F�V���]Qӏ�m*z��M�!
��;ao������^�&޼�\�8h*���F��]C
 К�	wq����sB0�?K�,���͔5i�jT2��c���m�ԙ��*nBx�s<�~�̪��Ĳ�Fic�]o�wS�}���Q"�`���u4����G����#��5�3�Oi�=��� ^̖a��[��'��?:I�դ�K�i Z�v����$w���ԡhw�,I/�e��ٞ�:z��	�2[]�Q
�q��	�h�抖P��@�Wx]DL\�q<����p�ǂ�kͥ�L.[��(���XK�� ((YFp/�z�+����E����͈�h2�N��21��#�ʽ�������������3�.9�0qu"WF���^xgT𚳥Y����t6*�vT5
����GPP�������!.�lQ��Y?am�A����������=�n�aP�ΪO��vu�"H��M�'&7l��u���j��!m��x��{V9t{���z�;��M�E���C�u�R!�	 �E�`�(3wgzy���N������Y[ÅQ:B!��I��#v1��-0�V"�H"Yid]��ru�Ep�M����b�D+��<��*3����I�r�!8,��#�'%2I��'�4e�ظ�x���Y�v`���)�Z�b�h�����!�7D��t�d;�`y��ާ����70&*�
���x�&YO7���|��4�+޽�~V �/��L:��+�sXv�z�Nn)~"��s���Û�]R���9v�D9� X��YD���A ��"k~0�+�q(�Z�0��\�q�ųد�ƪя���ƛ�6����*�*D�ƽa?wW�����!�9tS�^/J �	���ۑL�Sc-Ћ���,d���q��.�AjHK����M�����5��5�	'��C�-�
�8C�Y�W$2IH�`@�bG0?h<���K��T�ha�6҆��7@:���|��W��"��䴽��?cg'�+R��<Ay��2�%�,��Or'KL�U�ۑ��o4�n�x)������<�ڒ���E�E�rţD�B��ع�B�5��g��e���!����P��
\�t�d��S����ᆎ�i��ˬA-Q(��Fg3���6۬_��HT�5bڙ?X�~I�dm:V,\�/����W;@��Ji=)#I���t�_M7�KL�d�8/���Z=
c�;��gx���׵���bm3��S�m�0�vW�9$��1XTp���������P��f̿������P0�?����3�9��j������KV}(��/%gvmDV!H�� ��U1[�޼�;zP��oy�Z�w�t���E�i�d�i�t��y	�ڽ�K��뙤��K�L`���4��g�%vP;���&`(%�fA>��&�=��.U��'"��0Z���٬GR��^����$Ir��8�EPiGn���(tV���k��?�Fv���A�Ǚ%�i�U|��F�]*4md��>td� $����öR��e�$u[=Y�bM$-����s
�o��Y��`����0?�w�;�il�0c�y-��X(��!0���<5������k�B��t��p���꺦�`��ڬ�^R䛔���_��i�o-,X{�/�D0l�Ke�v�,��/'�0D7v�����/����7�vOq�%��'�$Pq����>|ɋ��@�!��ub3�X�60��*�H%��>q,����J���&���˚O�+@���7�����O��Q�U��qE��N��h?��	�ʜ��>r��<p7����n����#��:׷�s�|����e��r/�I����)������yo^��%޹p7��~<iMi����AB��ޘ�
��e �˟�^.d��0ro*�!���3k�YS��zQ�4#�m�ݰ/�N�j�rJ���~��%8ތ�x�bO2Bi]bI,�7|[�Î���V��D:�-D,���:�<5*��Q��ǎ���@\�wd�@���ٽ)f`Z"�����uJN��w�y(G��������|������!��#��X�i� ��3vJ��������׵RD�T�i$���
nz�>F%�4�)c0����6��v�_���uP�¬ӽ�z������F��0�� #96��&w�x�>�;>�2�üsL��q1�������@�C����\{U�\E���=f$VK\I'h���xl4�o��04�^��h\�\��f3��D�W�t����ہՙ��E�ղb��>�z�c6�Ŕ���Y�J}
�r�c���8!O�k~{1�40� s}��M�E�A���9���M!�~9p�+]*�&}�]�Wq�����H�$Gx�}~�9ϰ��R�dQS�]BH�L@~����f����l������������{�P�
�PދC���%�{}s�j�v����>�zS��6���N�}y��at��GxW��k��(u�!n,�]�������s�R�~W��J�hw�ցL��K�v��w'|��1��h��T0�n�dO�����m|���v�WH=6֑^�Zޱ���|Z��#k�(�a�.�_�6���֝/��T��ʲ����&��#/*���2 d���׆�1O��@���ע�V~����)�����L�5�s���H'��T&����V�[���E�u��D���X5yy���4��f�M|v,��w��-�.�S��5�ݧ<��/uqg�<�CS��)�d������b��
3x�N�X��=߅�'*����HH�3��.<ڊϧa�+���`�2��+���CӠنnn{�4ߪ���*|ʟ�L��;�1@�Y�ѝ%�p�����@ ��_أ��P*ȥ��ᑽ�t�����ʲ�?���S�x�h���p?��`u
�+��s�a�}@�O��EVH�'7�V�ȯ�s���eP�@�y�|ћ f��y�=R6��&�'�D����ͩ����<`�h��΢�[�7�D�8��*Ƀ��k�8�y�7>��ڨ������}�-oe�Z�̞ϛ��,��Z�CٵNp���/�\Gi5�j �޺Ʌ:�������&��j.T�2���H�)�.��� ���	ƻ.+�_����b�m�q�,�K[w�R=�Is_T�8$2����դ�<���f�⯰�_D@�<�`��zu��4��4�q�:�q�i��[��Z�,����_�K��7��*ĝ��p�������j/���)_�c]�J���I
�H�ͱ`��;p���()�6�+�~�S���e���b�En p�{��U}χ���b�Y�Gv�(�3�`�ď:���O��$�n�%q��!��]�[�#һ��fzrI\G����F���W�p�~;:��n��X�|)�����F���V���Q���{Q�,z�g'�i(q[���`,�٭;�+����M�`�o�1H�O��E�Q��nN}���-��0�0�1q�U�Ul��^;{'5y].MG�&a��(_�i�=9@e�)R��W�>���Q������2�-'�����׳W�n�CK��z ����,��v��+N[���< ����:�Vt	PR����C��^�e��3M��Z�Ifc`nnP�.5�#"�}]�E�*2 DA12� W�]�#����w�f$0I�>oxi!M)H�AoA�i�z.���_�� ��7Z��>)m7��5�c0���n�}[w��݁s}x��Z�);��:�i	{İG�c�#����ٳ��73�s*n��L���s�?������V@����F�-J�}�pw�s��X_U�r�RPC��[e��dV���x�z���Vz�G�V+�* z'����[��#��"��x�6��� ������/G!��F��>Խ���������z��TO�a�2u6Hh�f:n_��\��i㰡�/��s��e4�*�x�'���.�A@m�R���ɂ����G�U�.��x��t,@��Lђ#fn$��5[[�Q4�
E��i�|pius���_^n4HuA�����b��1R]5�b.B0�=�<I� gE��?Q�1ZD�[��W��g߰k�p	/�'��a����v��f�!�44S�1^��;
�馠�"�b� Z��5b
�Y���Ps����mG]��Q!���CR:.J�It�36�R���z���"}Q*�j�[j�d3nfd�L�~�Q��8��K�����<�w5�H�.>�a7H
2@�3�<�Z��T�Zn~��'5<�Vu*Qw�Vm����&�yZ��TD]�B�$��^I��`ck�9�F2�}��ϟ�.3j�������%U��0CS�f���-�������Z�	H�Ca@x����s��/N�s��G\bכ,i��"q �)}�����	�w�ColE�'��J�}�}�ɤ�2��o-9�0*�g %O���x���U����ی.G�dM)�<mJ?{��l.z^�c�>IIc��$	ԣ�.څ`w��,��M��m=	@B�F����l;��s1;���=>��e�c{�`��&��aM�8Я�����iX�0���HL��,I���bCu�o�	Ѐ��W��c�G|�oҵkl�rPlʑ|Go�6Y�AC�%CY�+�|��#}hQ��x�<��em����G���Tj.2c{E�6x��)s
I���S�$I�߿�fD�m���E��5�EjSe�W�7����R���ը��|������wr`ÍC~X�_?����<���LT3#�	����B�.������H���������6�BkКct��N���Q����Q'\F�M�b��!G-]*Y�����H	�M܇q��i�n��H�����-��i�r��:=�"��#�X��3�3Bb�e5ʫ�8��3��6	BDn��_��v� `:D���R�y~�����m?E�%o4��F�.2ъ�}ZO�=�aF	�l?�d��p�~}!Ἀ�^8�#@�P,����pw<Ҷ$����Gg
AqFG8 ▙
cN�T�!S��'�q�¸_��mi�ʱ���(��<�����p�TZ��S[
� ܧ��=g���U���ۜAb��F%�"����[��5+(�-}z�u9U	�<=�c��|�7l�����̪(�G�fw`X��+{�0����I]Ri�m���ό�`��z%���7F6Z_��"�5�G�����a9����~���rt����O#��4�u�b�9yǙ�������@�
D�� �L��XH=|��Y�L~���<���PN�����:�2�y�[���,_B��nT�/ ɍ˧��g�^��Ъ�ɖλ~go��6�^6�9I�d#g�5PGj&C1�V�Ď�]�X�� ��Ѭ�+3���P{�t�V6v�*f�A�r4ز)����a��^�wr��Hr���ċ�X�Q ԓ�)�N�=�Θ$�̜�3��Ky[`�o�Wۛ�=��]\C���Đ�Q�;�Ɍ�0�Z�uf��� '���%�"�ly2˿�3�&�K���̙�8�(�0Vq�gW��l�)���R���f��E�C.��<;�SB3��O�h!��16	�fr����2��I���s�ζ�Q{��x��5A�ͫq�(��@�,�. ����T��߆��B�㰧��r��2d���-m�WL�'�ao����5���bZ^Y�!y�"b&mM�{��_w禞Y1y��4'���I����:�IwV�%�ɰNI7f
��ƭ�q���dn-Yؔ}�2�Q���n�jw�/��x,�u�;��At�YoN8hn�
��tQ��)���ݭ��V�]�?�~��k �Aʱ�A�f`����Re��/�F|$��b�ؼ.�$Gp���'R	_�y�J��g�h]
��UqG��ܖ9��&�X�&�����5a�t3B�� Im3���sM�zq���1u�D���d��ʮ�
��t&���-G֮K#���ǥ$y*��QXM��dI�p-&�:q{6�J~)$��$��ʋe�)��:�J����ѱB�m%b#I9�R�l�d�L�m�4�.���J-^hMh��z���IN�����Ƙ���=�/�e�Pa�JF��^t�5��9ꉘ?H.6|CMO�0�40�}��l�P�؀L���?�Nk!�(U��0��x ։���N� ������ ��x�̡�>�7Jz�o?���+�IA����	��<xR?߽2�鳞�`�ᨲH�T�dBm�b-X`�˵�娇��'��G�6�}*^][��j��P7�9�{�?<�뼩�F6��K`���`�4M�w��S���{��-V``Z:8��s������p�/#�����s4�0Z�R@�%f(�ӧB�"x��̔��㢏��2�����3��,��pƅ���!I�If1�t�١�-f���I��>o�����C<�՟�6Й<SوZ�t3�'S��tl�wq0�	���zn�����~����M�?�ޡ�P&m��p�/)*�s�3��a��U6N����ܯOX���)�B�s�EA����5�>5�����u4	kB4�M��.%�����"aP�½�9H���ܙ�����*2��;<nXђ��X(D("��@6����w40q-J�w�`��|�.�B��V@T�&����>�sb��[�.��$;9�GIT=��M$h*Ktk2�CYa�#�fZ���'�)��:$��v�������g�%�R~��D<���K�Ԑ`�T�����YH2+�R��	Hu/�8��Gܜ>����e������2�DhhQ`�"u��*�:�X��!O%O�m�d��ଓ��\��߱A9��eo��I��I�d�:���N0����&I��T`���
Nt~2���k��Ƈ���."W�+��YאE���:��G0�Y�i��;c�I.�C0 d�i}ijb�k�$�cU+��|X�X��F�U�u�V���Iuϭ-���Qw�u�Z:}s��:j���dM���tI��1����6ņ�@;dIǕ
�;
�NTż����_CH�oZ��3��(���xD�g�|Aq\�a���ꈖ+�l/6s���i�2��H8ӽ����lE�Mw�ew�֚�U�:o�]�H�E;��+��[����,�2��0�"x���bZD஗U��2@V͕vOy>0�L\I:}�輨��7�8�;�A]��gL�8��r���9�'ݍ�oG Jx����ʚMxi���|ͫ8���}�g�ѳfB1R�b�\�4kp�n�������V�H�� ���^�b��G�wd� ���/{�f��1�W��6Ox|"J!��1����W���G�\��!�������@��%���A�&�����oH�U�����_��ʨ�#㰶U�V%&i8���%*]��,N���	f.P�Z�=j�l�&"Um�y-����q��������� މ�h��Ә�>�æU?������5����s�H���m�i���5�/1o���O[-�sa�{~�Ҩ�.���j��Ik^���oo���/l��7����_�a0Ϗ�K�PNyc�$���x ���$q�lz2�rb��0��S��������Tܥ|�c���q"v�6��4 M�>�z�s�I��V��J��`�Z�w�������
z, ���hf�'�x��H1����><���V)R	�#�*z�T\����[��4�����ߌ^�E���3[�m�mI���%v���ڊgOO�C��:�ܨT���rзT�-ح:I�+�G��L�*2��QY�@ !����
$����rI@������C7G4q��w�f�Ժ$�'&�pb��!n��@���g� 8�S˽�'i�p�x
���N@H&)��0�_k:��O.�h�o�`<��v�.�?Vf���*��6Q�����S�.��y���7NX�ׇ���o?�e�����V�� �>�zmA�������*<�*�Hxm
'*YaqO����S�ѱ�Ú�_"}r����w�L�Fu\Ƨ.̣�P�	s7l��x����k�y=J��N� ���&3~4��yE���|7��5s�*�t�80Qx%5�@(0��go�M��=.
:J�f�ȡ�v��-X�ۏQa	���kWz5U�jĿ&���C2��a�[��e���*�鲢�ϣI�M�$�ʘ�Z{������{�� ��
��7	�;�M���h�a���Gs�L"P�������g��$Jp�5�ZY��ݮ�S�r���5w;�k��pr�a�pˣ�����:EbK I �����7�2�T�P����k.N�S���X�ɜY#���7����$�63� �mj�g�C1N,0�Id+�M
G*�k˰p�Xߥ�a�P���M�� AQ��$ϩ,Q[�K\+�UP�,�|5�UxMJ��o��C��FBt9�1�9�b�Ȉ8%�'�"�ǡ����C'�-`�":-���Go`�0U}D�0�-�
Ĭ����~��gz\dV��x�CQ��h�	J�殤����^��кC#�`7B8�-=1Ɵlx�`~}�r tv�j�%�L��`�IUQ뜞�%�,:
|b�����b�,�b�9��v�K��U '*������2�'�sV������E7()���o��g�<٩���8�ޥ�\t;�-+d�d@K!�;΀�H��S�!X9��w��S��v����%���-vRF}��~�!�?�to>���j���n��$k����8+�O�E�0�x.�� !e��D�7f�m0Y��7�%K�7�C��=��0N��\�����W�)5� ��$Ƽsr�L�C�Eg�e.�G�M��~y@�E�s��&� �����p�5�'��$ ���J�����P��sm�ii�9F�k�����vh��Ix(@��HYLD��	�B�(�\�}��������O^��O�Bf�G�^�,��f�zn���ҡ]7�U���8dXNe{�ak<X�Є0
�=z�_^�������>3tΩۉ�O��* �ԅi���1�S�L����#�F(�����frא�}$�)���3�C|��]�hL�朂�>�y{�$�̽n��x��r�N=�Y�7b�����Ԥa(a�r:�"�s�`�QD��0�~�֍����k��k�Bi�����.��.u��_r�ú�3�X�9��kWh��&��+��*�c�˨��-qs��c�?tQc(dq��h�9'�I���`6@�@m�����.���:r|�)�kt��n�O��X�w�NR��l����]�5�0LI9�����9s��������=F�l���)��}�w�҂�S�:I��%�dsH*�^�9ug��`��{X �Y��`��u���d�[�2�6s��u�Y6ȋn�k�� ���;b��u��Nz��ׇ�)��ӑ�=��+�m�3��k �74��F��Õl���{W%Tcu���t}���mx�aG��� )����Wv^|\�8`"�ۀr�:G�:�Vڂd�Dw쏔J�ٌo2��z�t4<3����.=�D)�G!-�JG"�6�0��7��3�b(V<��61ֵy��N�Z�����kP�%C���W`$�v���{���Ҍ����_�oJ/����S$���mz>�!!/�7��-a9�C�kMi>E+��86S<��<��� v�8�`����*Rn��i+y��۩O�&o�-��^�fr�d���B�����q�<7'YHt �ݷhN�|M)���O *ڊ����Bn��h��	�o{��+~_���&�砹69���2�������9��9���fQv~a�����zTa{%�Q1����:�t�8_ݏ[��@��������OQ��_�����I�����/j�B��1/cg�8��}��x�V+q�����a
@� a{j�z8�h�4@�n��LF�aSg~,�Uv�o,(z��E�W����Wm�]������y4�v�_����p?��IA�(|V�9����߅�e��P������ufI�ɰ����uSԵ�XB�9�O���8zV�Ўk/y��� @'x�a���0�}A־�"�	#QH�vn:����i ���=/qN��/��J��-%B%:a^c���t��)��]%0��D�T1LܸGwj*��{�@��gjV�䀓�d,��o��`��"�����w��hYg��r�����c�Yi�Dﳼ!���[7Ӷ~���t��p���}yj��TK~����\�L�x"aM�'wG��=�K*�m��a�I��;P�u�+�ȅMI0c��H����tD^S�W�<T���%�<�T��3������6�`��'PN�`��RH� �8�RNz2�0��Z����NL�`u �Ub����L�M�,T�W峪�@$m�@U株P��T�R�F��;�H����>A��z��,���Y;Y�$ԢNiմ�P`8�ᥢO�/Vt����X���n�d	N/�/�����������:0�i�'m~��_C��%�K��)\�9��+iW�5	}(��s/��V����P�����%�D.��=�^2��քb��\1x�ϓ"�'#z����Z[w��K�����xw�R���!��m�C�h�0n]0dy%~�~�Y�228sh�����Fiԑ�u^*�d��י{|�e��Y ����;VȚo�{�~��լ�}G60܉��6*%�P��"s�Yd��+TjP{[���h�����BPW�3S�s��|j�XXH�[���6#���{?d�@��7��o"Vl�ҥ��,���q�.�ur�\0;k�Qh]t���Ɛ\@�E��c`yA�_�Ėu���a4$I�ׇb�4b�a���<�N��c�����UğH��K�Jk�{�4_
4��h����p�ŎZ\c�\�nwm���#��f�(m$̮��хu��Q$�v��73{��)rE.��_�;���vT��U8��\��o|~�f^7c*�7��}I��kj{u7gzf��ɼ�a��s�`Т�eI�} (��\�o)���5V�>�-������uLk�$�AKpm6�\[&	��<J#�@B0��S[=� �Í}�ה�Ϗz�����S��\Q{���Τ��u �t��ox�"{�2��t��������&�����2R����<�ѽf�ҝ��w��k"!�R�s.aūvޓU�J�q?ߋ�R��V�Ae���[GQß��Pz&��̓߆Y���7���v��#��ʴa9��T��D-lFc�p$��'����B�˚ǖj>(��CfIyU�����;RH�|F?�>@|]@�Ÿ��F�QoHT�4��ӿ]��B�	�{A���p3(�F�����S�6��ClG�vh�I��9��̣��\o��Q��N70��� ~g�hXh^q��1�^D�n#Br�����d���[��l.�OJ��=�h.���te��*�`E�:���q�A7����&��;� ����P�
���""��O�u	S�0/<H�����y���C�S� ��Ypy��f��	D�����G��׷��pg��\>#�&j�+Z�S�l*SZa��s-�x҇$ж[Hi�8�̒��.�	�f���Q��|ʬ��"e~֨�K+ű��)�
N�K���M�"H�Y�e�z|����gm�K:�a��v8�";9L�S���J7����G 	1���q�.݉?�A�C�u�Ǡ��Ul;2Xs�'?�R��q+$o�������1՚"��"���kn�J2�ީ+H�X_�I�VbaFM70��w����4@���H˫���P`��$�d@��`������f%���ha��o����0���I���#�-Y�g�*����VK����L-k��#}�i5�0��*��!����z\�{�VW��1|+��A'n{_�u�ߺ�0����E��qV��c,��2�添�9��3<�2��P�s�T-꒯�	�p��W"2�������c��~�b� ��h=дo��`Y  _^���ߗ��M�
,�q &'�	��߃;6�5C��p��^�xt6�(��[��[�(>��V�=��l~�X#�?ɍb ���߈)���RˎЪs�`�z��k<��o�{��Yh3ϟ����g���+����`���Ы�K���iV���w�E�' �&���zq�m�h���Q4 ��m��YP�J��Q�&_O�7�g����aʌ΁�y��@����N�r�s,gd�I�-10�t�t[.H�sQ�l*�B���G���K��|�B����ʕ�����AW��6�|G�8s�g��QՀ�?De��c'hK����rCr��tg��q�����x�ځW�("n`��7�؃J�-RpR�N����1d:��I�=]�����䃾Qg4�Q�����L��w�0�S�h'q���T�� �i��Nw<����1�����(��}bB��PsŌ>F'���:�y�����44M�pT~TYV�J�.b��>����[K�����j��Gy ʰ�YWC��;+ZNË��3��.�9
�*S��@��D$ԃ�3!!�ʳ���շ���_P^�[�Pvo2流9�M=>O�}�3v��/��:!v"_�Qe��d[�m	��/R�{��i~jw,Y�(K�@F����p��(��ǿAiN���\r��۔�Y�r���1t�����jb�ܥa�Z��;�أ���e�;ٍ�_`i'{2
o�V&�~E��ɧ�A;��������pz̴�	�э�������m#P	����Y����$�~�%���PoO|Q/0N���S��mj���_�k�v��IG����C��lkh'�G�8ㅚ�qP��_�V0s��#L����UF���h��q\�`,ƹJ�%��-�嚔���'���5��6���d�G��>`�+��"�!Bm^�a�%/Q[A+��|v�v��ͬB@l�AT��s�S�����mf�[�\*>s��ӟ�#�
w��*�ꍛUY |ߢ��V��¨[��c��:��%�/�zҞ#�f�	��n�Ϙ�\���'Q��0�P�\u��Y
��^CH�f�k�?���svG%�,G�.F%?�ⰻl�Q?C�kc �h�j�%Q�u��p���{�j�9,��
|9�i��B�� ����Ze��'c֊k��s�5\����_V�����eضѭ�ژ����P
un�'�?>�������Ŗ	-�fOB{J"w?h�ӣ���.שBL�*S!<�b6�_$
v��/�P>1p*<~�3�$+�}I^�@Ĝ�'�=�0En�GhǕ�@�Eq�Ĵ� �?�&��/�ߛ6U[lv	z��R���;\�V9���a!#}
�C;��E�3���$�����K�+�J�[��:[#��FHsȠ;)�o�ǒ��fJ��P�v��"K�%lΜ�AjINN�/� �`qS�鲢pe����A�',\V��i`+�d"m��>���S;ڴ��f���#c��e�!����E*! ���#8��<����ʋ8I{в�������>/�L�o�j�l�b�ck&��v�=yBCJ��C�5M��U��5_�뀣�����`5:��zo�2�\2{�Z/Jj [�}-DЎ�X/FX2
��{��~�<. ��[F
��I�z[�)�� ����+����Y3����k�y���f�_0Q���>����^�R�38-W�
R(9����5VFF�`@���Y��쑁r6jņ���sN�*��|����4L�S<�hd�1R?9�R�C����a\mՔ9�O������]�:8}˒ּ������3��i/L���eE�J�˰y�M^4��VQb�{�9�i�g��[�G�aaЈ(��q`M��-^���UE��~��1��ʤuw9\����i(��;d��*TZL�w�ݐ��2&�Wǘ����Ωf�{vؾfb���J��U�3� �ד˵��K�{�!��G�wJ�	}��i�z$?��� Fi[�aK��u��K�l`�	�<9;"���'�.MK��S샷?���'�����Sl������<0����'�j�۲��� ��z:�mR�y��(ڷF��w��(:��≾�8���!q#���p�I�w/8��'3U�?��r2V�I�:�����_�x�C&�)'����fv�2���s���=�&v>na*s�)���?�i�p��)����	���7��L���e�	(���P�i���~�lo#�P" ��udO���I��	�^I�2i5�����Kt��f����f���-s�Sk;����v��$(ɠV� �Ќ�s���ӌPM^��A�������L�l�9(���a��^QRqG�#�Įcp�d ��K�B8�
'�	c�ǶG!�g{� ��')1�v󰁚#�}�0���m+�f���z��YVX
]j����z���s��9A���/�*�kkuQ��-�"2DE+AXv DѻZ�_��L�^	?P�MgE���u�}Y������r]ĭ2#��:���qǉ�1�Ԋ�w!�i��?l�$Mto���ɷ��=Ÿ�66
q!���~�VO��)V����Q�]_}��q�`�c�GW�����uO���.|��Q�z�*�S+�$�������-(S��B(�pe(Q_�n��7�����`b ���;$�pl�мf|ԧ�m�q���$�l\vV�Mtɸu���x6�/	��ɝ�%���'Nhமhvm��v�rS�N�װ?���D���6{~��X|�R�Z�|Kb���fiM������|�;��=mM\]��o\�_&�p���E-�5��p�����׃j���҈(�0�K��]+�,� ��r�f匬	��Ӆf�����&�VM4�̩�(���$U�������T�OJe��L�&op�������_��u��, ��<�=/��v�;ϸNV7�r�n�d�g��n+�V��ox��ɈN�9�7���:�>�p�l��ڟR��:c0�f�&�xu'��UF4y���>Κ=R�nY��!.+�Nl����^�pC���X�&6\_E��GT�Å?71[��������1�L�D�W��AKK ��<L�\�Y?{��*@���'���{�da�H�$���굲�o־�!
G0�l�:0�w���J&�p
�������ו�@��
V_�v+�O	���ү�����O�{M[U��e� Ū�lS�Jw�*����:`(�\�"'�	�r�t�y�*�zyGP�W��$�p�0ÿQ��!K�|����&ͬ�Pʲ��]��G�A­՜�V�\D�=��@�x���u�%[^˹	�)<ӳ��|bKp�r&g��8�H|G�9�	�)\q~a�3���5��9�ʽ;������wa���X�Z�@s���O�c�����d��;�8�j<�h|�sݚ,�<����9<w��L��}���6��"���2�z����HA�`���1���[�������#}����Xz��� Ա�@
<+� Y��(�B�y���7xhf�ϙ�]Ly�v�(z�Y�x����SM�m."�캣б����F�ez �XI����]w~y@��
�S>-��P;"�ev�:� ��DC�.+[��>���ʞ�;�Tf�����f�}��2��x���qK�E�!W�C*^�L=fit��إ��N*dDh�d*��4qctrB�12�z��t�m�_�X��<Po��A�X�;��Yz*e���v�j��@y��ƿ��d�D�K�+f�]���!���S���'��<�����ӝݴ���D�f�p7|_3����b��V��O��5�z�Eֈ�G���ZD���ů���3*xC�a%*v�6L�T�z���\p�8���|�0d���c	�.���g����=�������TE�Cu��L��0?'5�Sa7��w�D}��b'�y�O�&	5R�d�i�|�Lv����iDaqk4�qI
Z8�d�cE�����&7�F�]�Z)�1�}I�̐��B�P�2Q"*kY�P�_Y?�1aj�u� {��h�	2�9ǧe�d�ry�?��g��E�,m��R�z�Էk��E,-`��U�� �cu�����C@����(�J�Z����z�jn�.L�]� ;�yx&�	E��d}�a����%`%<p�-��jbT�J!^��<��ֻjo��93R������ ��~�Qs�D/M�яK5���ih�p�b��v�x�ˌkg�a�p�Q�����$L��k�`�"H}�жY�U�����n�Q�������\w��s�5d����'��؏%ٰF��$�j0,W�[�R�r,mZ��@�@w ��pl�&�$��_��RD����������{U��%]��x~E+�ax6��+��d�>8D� |o�~QV����*���Տjs�����HV4�d��7{�G�q>��Nfr����?�E���E o����%�w��J����0r{�XM�(X��ͳ�5�*J'�d���%��1�X&�H�=��h�{hk0� ��ށ;�p��٫K�|��8V��\��8,�~\�5T���@2,d�!��X�ve�IL��B�2j�j��,�)Z��.H�d�!�����D",G��h��(d����t Q(�N�|2��W��a"{tj%�7��\��X��G�#���3��U"�Ln� ��h��A���k(^�o��_�h��]4pU� �Gtr�M��hy�m��T2���vK�w����X�nR�N3��6$��Q��rWJ�z�����]R�����l|�KF�Em���y�=�gQ,�$��{�R.L1����:za���t��=)�Q�����E�;�L��ɸ;�K�s�:��~k	QYڡ��Q9�c�o�$���$��6����Sj���G�d���zpO�u%�X�G�V�<�����w�o��@T9t���S�tr�O�Z��#���S�p��.�NŘ���o�ht�s�Č�q'yB}5�eٌ>�peU�=��mk�+�ۑ�����Mi���+�r��n�;,D�X��"#E�y�(�y��z��	覀��Qq��j��PL������k��ë���0:Y\���h>������ 	�����ᶍs�R����k~z	��|��b(]� 뿣re(�u�1�b��Bjl̓k�rBY0�������XS=��|г��H#,������^�*�.Q)���Ao�9V��mC?���S%�k�3M�,�������^8�J�	�kTE`�"v{��8���.�q�fI��Q�,t7�C<`�y���ހ�%y(��Xc���lsz�~�g5ē��!���������g"	���8��8uJ��
�?�@詶d����.t��ej�~����	c&��oa�Y�_�%3ggteJH���v��#$�4��/�n�OQA� ͪ��Q?ʐLI~#�`X���r�!u���tт[kC�
���*5¥�s8�o�DˣW�7$��f��pFM���T��$����@[���&�yx�,t$�e�3j5]v�W�i.%T�o�����[� �Rd��m�X-5y��&@Kh�	_h{~�?F�����l<������K�ĝ����J�<��h�M(�/?9(n�����R)���?LM����Sk:�`4�%���������5����F־JԎ,����=t�Q�g<Y�`B�5]R�$�4`00�N�ge��-j�E���]k.���-�?�%s� ��HI8�i8����?��|��CA1ƒtF5�,ׅ�X�Y{IAk>�v�ϑ8���Q3$�W6����MSt���"8�xʯFK�Xҿ�N��6������e
,\�i�B��OV),�ȢM� Ϩ�⼃'�8�3hH��f|���Wv��gz���9~�6�.���N ݲ�1�a����3����e��(p͠,��4}=�Y�Ң
Ĉ��$=4:o��0�Ȁ�q؛爐g�V��p��.�ZUo/X���$"Y[UU��R����"tfЫ��o��Q
N�.
6�U�R���ǹ߬w'��-�y�/�,(����2��$������W�[_R�3/m�b>|O�eR�1�a��#Й=�1�1n�Ն&�#W��q�?�+�݄����k�si#r��PM'�
/�_)��N6��XN�Mn���宆rژ�܆rD��h��1�fS�`�`]L�.*���u;�QFJ&��.�5�'=���#�ѐP��Ut�;��=e%���L�����L�p�i�rӡ��M�-c���J�i*���d欓�(�G��}�^���h���T�E�!Ȁ` q����\>�g1�tE���2r�7���@�:r�P3��|J�z�����_+>cA�{>y�W�> ����xH�� �����v�=�@��LL����*�Q��.�3��	���OY��Yw�11�fq�ړ�4��s����,�󾫐��w�ڙ$p���^A�^���΄c5779�N?A,v�eդ���_�=��E�W�,�|�g���y��+�Dg(R�Ւ�7,i�|]_9oo^�t�X�+��b��pG�gA�����JA��ZTW��q6s͉����}��\���۴4S;7ڄ#P��W �ܕa�^�;څtP�2���;����cv�h(R�������(żb�_�츼!�^3.:�x�-�+��)��db�ޯ+Wa'�ύ�0���33 �t��
g����e��wP�$���"�<���c���ʲ��oS]l�(��M.���	y�dg�5n�Y����J~�1qA`�@h_��-ǽ-.�1�Ѽ���䒺�����jYėݞ.� �����趬��-(Ǝ����X��A�ǁ��8�WJ���a����J�t�1�`)�v)����9��b/��KMM`*�-���<�5��'�b���]��4�+�(�q�:���}*sAEn8�"���I�487�zD#�@��Q�(��(���-9�{��t2c�[�x����E`6��I�$t�<���|H�Yʥ���Gy�4�:^�	1v�raT+�	ӗ�_�\�Q^�{`XuA���o�L_���c���(��cm���{:Oj�hW6N�߽��Us	јb7�F�֋��.0�xY1םFl-V6�E�ϐ@=���&1��� ܗ��%
���'^��Z�)�u�CR��gď��U��EΒC�/�X�z e�����ˇ��[r�Cy��CФ���yZ�s�i�_���9|{!�Ip�lt9�h��O7���LrQ�^�,��f5����L�,WXs+�x�z �^F�D_I=���N�@�!�n�j�f�\	����+H��R2K����\��eFբ�g\
�9���q+��+,>9&�����Z�՞�@&Zc }���m܋�$YuHڐDl��k,�2}�9�ܿC0;�v�i��f�-ՓB~?}6�;p����(6Ib2w�\3�P]H�q�"թ���u!8�B��Y�<�^��Z_�X�=^�cq̃/�l`�рYD�\�kʈ��|�TrŦr������Ժ�#J�ޒ�kf����R���HE��˻:�z�.�Ӯ��Qɗx�Q��FŲ(g����/�ƒ.���@;s���Zh&#�`x| ��٬v�q�6}�R�IP$��Ŗ�\�k|���h��|�b�u�^�"�8�?}Y5����<�gAP�3�_�jV4S��eޮ���E,]b/�ߺ3����}��
���@�����Q�Hx���6	p�$	��W�p�㉚�Sy���{�4���=�4�7�%�b�fI� �kN@#O���F(x���7�;�`�ֺh-m���_��u�(~r�T)g!�	/Q��>�sj����܏�|�U�5��u�Rr�&!]N��.Rd\�é(i�d\�K���O��V1�/�kc6��.�+7ԩȺX=��?"�c'U�s��3'7�N�B͝��1�"ͪ�*�����hd>	�.M`zDUY�N��/��ߟe��Љ]^r_<�#45��vYt���]� 5��|���%���X��8[h��k�W�M�<�+�����/6[zG\�LҏG�7̣*U��=����8S��(TT˴D3�BY��J�P���a�ܬ�Q;�C��0V���U�����\l�l��O�Ʊ⭔1�(�ճ����F59��9=�sC�ާ{nD��Ze)�#r�.TIq`�C�f��B*Sx��E���O�&HB��:t�!��wT�M���?�Y��f$C'd�.b�n���b��pw��#\o��-�t)׋��|/�w�������}<�̍�XA�u����Nc(E�E��I�Gu�jY���C#4�K�5�]��_�L8�SLuǘ�%j�������IE���2���j�e�´�w�] �Ť�]2}�%t�:�{�*oO0�+y�`6�DU�.?�1��޹O�4���<�3�kLN�:�MCq����4��Һ'g_,4O[�'u��i�Xj�o�e^z��C���;���x��#�v��<�����`�\߈ڸ}�h�Ͳ�g��!�N���2O���{%����\�[J9�Vg2/�,�~��{�UKi�.������*�WK�H���������N�R�P��|�y��j���1N�&�8k�S!�����s��1Ԃ�L��N��;qaL5��$���(��k+�e-sT�B�9�EF��,�U�9��l�T�q�Gv|i03�&�ƲP)%z��Fh�]IP�z���AI~I�]-P+�	#߫Z���)S}�OͿ����vf������l*51;�ݏG����-�`���� �sw�Lk��]�j<N�(o���	��S�#�+@�С�o�p�������t����K�>pP�6s�[��i�\��7��^�p	v<�T ��K����L�$�=��_"!�+8h�.������Z}v�;V�rX�y�/OՐ_�|��NR;Y ���|d��	��M9c��0�Q �YC^-�H�	GN�[��h��B����0�`�E�Š9g�xY��X�qu�1[�����ś�t&�>)D!Ұ����po���G��9��j�f�m�Y�3[�	OB=�"���'|!�n����F��A(��������a�h+`������U�f\�4�����'����N�/�H5����v�˗_J�F��}wQ��i�#7R@7�"�\M!�CF�-����a��^ §����2�5�;�H������tg�͗���p�ֹ-��7L+�}#���@u���{yy�4+�{��E��O�F`UAբ��gT1CIU��A<M�\m)_qo�	�]G2�����j���?��qΏnA�^�tHD+U�ۄD#}wZ�vŗ*yC�����ݏ�ԝv{�hQ���% �|����1�>��dr'�8m�T+-�kN��)ָ�Y�rB�S`��c��8�� �A�M���f9=�xR�M4
�X�jS�	�U���y��ٱ�ޫG	J(�ЙWG���' 4�G--Y1M" &̷�d��1;X���1fd.YM�&�돒����v4czfS!�F2綎�����N��Tbs�E�<�FM��^g�%�M6w
A�N��(̴�hϘ�$a�J'j��
���q����3�&�h�A����<K�Y���u������m���'6���r ����D��\���$��c�^b���xJb�we+�ذ�ͤ�n�F��2�����V�gh97�� 9�h'ׁ�yP�O%f�?(��P�+K_N�����|�P�4����"���䮧�	FfNK����u0��:Y���՟��k�K,Tڠř�+Gq�$�=�m8n�R��1�{���K����V��������Q?
-�|���!'L������["��"*թ�yڱGC?ҳb���w���A{��a���g�Z�)Uϵ�l�a狁���Nвǂ�[<�)�[J�{�A���l��|�-.�
��8��4�� ͓(
x�J�f�����	۽\�`Ҽ�}�� �]�xT.�`5+��Ӣ����^�����	��̾��1RPs�ہ�V2	F���9��I2{-@�:�N����u�(�	=&12�#�+t �t*��5Jm7��Q��=c�b�T�0��+���!�)z@��s��*U��jveBU��J@$P*�S��X��x��5F��`=ξ3�2䵐_R�X��!��V���b1��c���z�_E����yq0��Ÿ3wc�����INB�
Խ}cl������;9�?� T��GG-y�=}����=y"y��A�<p�	�������x�5������M�0>�6^�qk>��v�)ݍ��[w��q���R^k��R�t;P�S�V��*���c��3)�	��I$��vġ+y��L+Ӿ��FJ�.��$�9�^m�s�Ɏ�@������D�p�T�����>����n�����S��H�6��ZH ,.�p����\mSt�! ٦�}"蒏���Z�y�N������Nk$��Ƃ"ޅ�{HQDm��OW�AH�'�p�;=��'2����B�;��l��_�)@��.�+b�7�gS$���s�F�:Q��˷
��{�ƳMQ��2�%�ube�hɄ�`�$��W�-\�t��מ#C՞�%��Zh[R��\����j���~@�adǭ1�1��艒uY�
|5kbĀb[�g�hM7�G��)�n�U��;q�Go^���¿C*��0�=�=b�U�T���IM��S��Dnd�Ge��a)\q�uw6��&.U��X�d.��a7ULs�QL@�ڃ����Y<R���\����5��$�W�_R�{��ޕ����G�0����Yt��3:�Z�qNh��Ay0���_ɖr��n���ݪ�I;`~��5ñ��ٺl�;_���y%�͏8X����I�Q��uh�����XG9g�x
d�452v�#�ٞ!�5"_5�K)6�Py���ˤ:����c1�#&��O�����9�H�i!T	O9��U��\�'�~Щ�!�1c>����G� ������ZuR�kw2��b&~���c����������4��q+ՠ?�.���3�'9 �DˬȎ�'6Rp�ko�V|�x�����a�v���y�� 2t��B�ٯ���Ȅ��m�@߳BI���c!ýq�������	��_Rٕ��,}D�m4R�'�)�!^2����4���R����T�D����G&R=�	b���0��,sd�"X�/?����{����=K��0
����a��?V��Ad>�/ 뇹t�q�����(��.M���VR�L�;�#�-��C4�ᢾ���z���)�I3��I]�9Z݇#� <�~�L;�:Wy�z��ÿ�ZZ~	��:��N��>\���1��{$�U���	�[��l�({X�%�A	+c�����P*���$X\O�!#�N|�0\���!��M· 
��u���:w�CU�[��zǶ��ʼu��K��ٟ؅P��DUTl�'���_�u��=TEId��˕>۸.3����|W���j�I����i|�%� /r�[Γ��7O�62;q�b��I��j;���F+�M���ikj ?���P*��Jp!�O��%��
�A�3��	��.������g��o{l��'A�c�޳� cI�r�W8$-������!g�
�z|��t����QE]�06��7�10�'?C>��.�3�>c�>vㅓ��Z�����HL���[7T��\�k e�p��mQ���?�&�lO���9$�[X,�d8��qi�����2�	r��1S�&���|��nb��%��f�+���}pH������-��=S1��Y�J��}�<�ēMʤs�})�i.��ݝ�}<��8&��io*���g�{���1�p�Or�h�g�f~k��m��yD��ɭ·��̅S�������L��C��I�T��e��"R@�e�6_����R�t>�5��WRa�>5A��L<�˰6<2_a>�1s@rag����-��B<X*�HV�����+*�C��
������D>��ҨC��4M��:�[�U|g�>
��s�K=��I����Q�:�O�?�Wq^��u��d1�݊X��4#���!��W\@��w�,�7񒄆n��â�^1�y����q��}]��].h)�3�[�ʯ&�<����˼A������%Iw�M!�)T�,m�#��``1�B\�>���@f�6K�U�8[��؆�#�~�|΃ך<u��\���w�#TKB,.�9�y��M��?�̸��1Ɨy�v?�j�H\I?�M�PC+�G��bs���!��R�f�Q� ���"�4�O�����/��[� ���-�99�q�DZ8/���~�������]^Z�N�_|��ˇ�Cf�H��M$9y����-�rv��8z��+��b
��`��6������u�Qt�������O���`�Oܼ�*��uй1�����#N��c��q[��"u�Hǈ��jvVg��#R lk`�i<��Gj	��5��Z��:��i�g뜣�k*�N�K�HxEk�7}I�l;~��o�l�xX���q��)���I�i<�	�n�N� �k�������w%��H7�En�<?���-�D�P6�����jbd�R�l�]�ԝ�:��u�֜.3���H��[ܼ���ǳ���E5�.T̯p#�
�3���mz� �ZEA]XrV/t:)|���,f�=JF~�'0V��fQ��ۼ�K�g�9�I�(́P�����Q�0� ��Gl~�+���ߍ"+�7���c`6�Z�S�N��'Yy�^�%Aݥ�-�8��--��)��3�;g�2 ��)lق�e�C3p�S&_.#7wD�roq�����7�A8�z�c6J(�LG��a`�@�>v�N��NGŽ��@lIa`&4em~�e����o�R�p���j<�B����%�ZW�Dj�GQ�|���T��)1g�%����_�@��p���x�������N�s������7&~犾�PፄE5�Sj�M��b��HA��Ѡ~{j��L��	�&n�m���ɗ:ǚ��ퟧ��S�e�o�C����ĥ����o������ 뢙�hH�.pj|���Ƅ���Ԧ��q��5����it���J��}w��ce��_u z���4)��J��(-���ۈlYo�Q������t��������R-�]�]��Y0[;�_��
��YI��B.�-�t��(@m��Z4���\�oiuR�Hw���]hb`�F~xj�ed��{ ������T���� xU$z6���|�P~v��=
i����awӜ�;{o��>@�{
��"�<.w`C�kV<��V.t�,ӟ"���#��0,.�Ҩk̾/�}�4��0��7��g"H`&x��=%=��>��PMlW�p���A���v1�E�z)JI�gy�8�#���l�`�Q�7�w�E�L~d1(��L0C��G4�	NXD�9����iy{�����zg���}8����I�6��,_0w���4�$�t���TX�1��8�� �f���ԊX JN��FX�6���>����b+z���}�X���{��ʔd�7��۸oA3C�嫸����,��i^ �P����2�#ݱD2n[�J>�x����n����L���4Г�x�2���5[�\�`�㼿�C�vӥ<3b�XqQ�oR+ڝ�X���ګ���P]�q4���Z��vB��Û�Twq�2��f�~|�%[w)4"�G��?/���!ث�����Q�Pm�;ߖ��0��l��F(J����O��,jg[�3�o�|�%�Z���q�F�8D�����z���"��V���6�ZR���;0r֨���@Ф�HI/�+�D�D��R����=�8�D}$қ0T�/,&�VSg�d_�����aPQ���f.�/b��Dc(�B̃�����߃��B�Aju!�o�(��G�,����c?)�M+spu*��_��G�t<��<�B��L�+_�A�U����;�`G�
_��ܛ%�
s
:��w���hl�j$I�����h���v:5��1�D���vȔ��V�y;�������=�\'�@��%�s*�%�fⰈ�EgT�b]R0��!�m���e��$��_B)q�?�Q���k^�HR��՝a�� ��Z蚓�{u�����+U���*��n�
�Ax���ϓaBjIh�\��h�N*�o��爐�|�غ)E�`!������[_ipaS��4gZ|	������70wt�������_�F��2o0�,n�z�H\����\j�����RbP%�2�SS��Y,T���2q�Tb���Z�>]���`!�?ɾ�&�Z�x���n'�p��9�W^�2�߫]����S�4�W]D�qG�S�d��n|�Y�� 4NAB�6a!,�i���T����S:�	.����F�)n�F�����G���Q�իϧ�Qx�L�9�*\���Ãz \��#S����	���O,������9��FY=׏ʨ�r)*<�@���(q�e�Xz1)�cS���3��I�m!�~�ę���-B�j�^� ɳ�D�NJ�?;ט�B_�C��Ut/���+f�og	��y�tL�9Sf��8���)r^A�Q���>p�y8Q~���\��ܨ�#Xq�V>�nx뼤v���v�A3�fiBz��^=�8y����8ռwq��a`
s���}�G��k`��Ѣ��ц�EiBʄt�}�����C0[��4;�:|=�A��e��I����ܝ���d���CL��&���a���5m���{�H$��ټ_ǑۣU���p�d�h������.��V�z�SЦfIe�Ep?�0a�.|����# �<-q������u�WY��ۚāBUF�()J@���&���ˁT�o�k;�{� b"�=�Kv�m���OP���e��>����˚�A��%O2)��K��o�7c5����l.��_�_$J�B.f�<�/���j_��"�.X\�k@�:l��D�lQe���6 "*�X�e�화n���K��8`ZD_B1�zr��\��PB��_~��s�]�p�W�2C������=��x��L��J�ƪ��]2�2�/�2{(.E^m/�	���k��=g�G���$����\J�I�d׫���t.�d�~��r����$'���- �ӎ��r[�h5�gQG?lЧ�X�f��!���.�;!���G�y��q����Y�W�bU�C����4���d�3<�פ�On��� �IB�ֵۣ�MO�sA�Ab�1���w�E����5�Ե�T�I#���奝W�4D�[!�OB������T��]o���]6�F������Va��Ť!�<�N!�<tN&>�r�z���A	�	_��%���	,e�!��.I_T�7\��/�L-�[E�+�4�w�\l+^:�j���
��y<��
iU]����Ż%;r����#RɩW���i�NX�MA <�KÔ�`���@��4���b�p�	�#Ҳ1�����qR��tgC�� eV$�M_�vQ�`�q���9ɀ��5X\X��Ҍqw�]�?F?���?}��!��K(�XOq���Y��6�/�%&�f��`��Q\�|�ߚ�+�,�Q�DG���s�[��u_x2ȉr�ph��5Ӓ۹�I�W��H=�E��C���kx��p`M�JQ�"���Y�������Nݢq�j���=�2��ߔ�qb��8�yӼ�7y<",�I'%�Q�8>��?�$\SU�up��!NN�~��ՙ|ہ�c��R�`��)�u�.L�ih%�)�z	TSts\�1)����­�]#���<���J�xmo��D� ���s���Z�e�Ⱥ��J3�'K������X�۸qGE���.n*bLZ���[�1W�z^���fR̞�w��������NQ��E�'����vb'k�WiЁ�(�wz�g�Œ��tu���7�2w �r����=��ӑc�"F��� ��M�He�w�Ia�����m����E�E�	Z������|�X���ð�d��lJ���hëc������l#�_ަsD��Lo�4����?z	F�6��Q����P͵Lt/ ����%	�	��^�% 
X5҂�IT5���|-㆕�_l��KE��uT3Pr�pn��(]5f��gr��K���L���8=��B���f�u�{��<��|ǃU�/_�( ��r�z�rZ]5�~H���U#jT04��k�S�w��9��\^)ƕ��Ջ���C��_�]Ck�~=�@�lх�=���dY���w|E�\D��n+�ܡ����k�o~�؍)4?4N�ss��SJ?< Qn��Ja���}J�烠B�U����W�3���9�?ځ�5�Ј���GJ7��q�* �&W$�5�~
4o� �������l�٩e	�
W�],#Ҍ�M���/��g�LM�"P\��!�D�W����Fq(����0���9g���&I�����w�����|Ad�x����@�m�)�ێ�8��H�?g�to�H&��f)�0S-c�y?p�Q8+��u�7��W�_�W�*�r����-H�,��|_��F6����FE��&2ӰM�Xla��q�ƊTMwCaKD5��u׹8�?�o�!��qʙ��Z��}f&��5�2���ho����e��+5�|�nٍ���B����`3�e&���[�
=%��|B��h���w{M�΁=��?zM����5��NnAb��&�Yys���a5�B�{Z=�L�U�:���%�6�5Hr��/ɯ��7��7A�x@	Qףݰ/K�RGB� CB{_e�5�E�q���T:��]�4h�����0�T�%}|Q�KVBu ���Fk" D \"�Q^6B�m�x�Yĝ�t�������2n/
��3�w��@�hl?G�)f��XA7(�7�t�IB�R����t�5G�9z�ѽ><n�@	�E�&Mv���D �����_9guL1�͊�F�wOB+q<o��	�F�Q���� �D�������V��N$|iU�4��֖%fԠME��i�ZDB��\=�ܶ�
-^�O�H=�j� W �l|��]�['�TF��n{�:h.���[x<Z�`��.Zi̭2���jUƦO�4���c=,�*�W_XH4҇u�=Ļ#"�G�笋�41V�x�2�`��o'x�<(.�g����6H�>pP�u�F�g�2�������z�;����Ld}�b�SE��)�;����x&TB���P	�ݎO�P2o����G�ΚR6s�oq�:�Z:'�Y�^V��2P�� U=F��p 6{>���� �����Y��S����M^��͖Mfڲ��xc{���rB���GG�a�Rk"�a��{�ehRL�N)��vF�J�'�������D�����79��y��ͨD�Tn���2�Oe�tN|H���C�!�$�lWծ��d�pT�A>G�@Z��������t(c���ZŶݷ!|�SKH�l&��`�^´l�ߌ����g��ǅ&���vF�ϴ�a{]��7d`.-�(&��4�����~%Y�:`�g�:���/�*���z�������1 7\OrW��9N�@����?l�!*��IG`����n .*q@WG�Vs�����$�'^Y� ܻ�\��G�m���8y�!�K _x�F)?��Gxú�9����0�J��=������YVfxҪ�k*��Ќ����'�e�`�[-�Ab���E�}7$�Hd�8���::�$�aq�$�M�w�5Жa�:�q��R9*~^�l�AF|燆P�s�-��\5��R�{�"C ?r���Oz������=1�7�	X���܉�P���͹v>\�����@�nn6����4P���3�2�裆���F��$}�Jl��Z���yy�W���j�6���M51��_�
�e��y�x�ʖn/:�x~\:��yW�m�JZ<r�=^u�������б��҉r����5
QK�'i����L8,����}d4�/M�#�����h���#�|yɜ��r�\���?7���>E�B���^N�3J��u!�Ίl�k�`�" �9���7u�Ǌ�^�b����E����յ�n��,mwX��m��ܒ�j�u��l<u�E��*�$��;&7��*X�'��V{;وTGx�S�g�]�HJ�
	���e1��py%�jౄ�y��9/7'􃍙F�(_�Z���:$k}g�a��8���L4�l��U�L�vc��-�id:��˯C�jТ"=n�Ȓ�o��͢#�y�6����t��.�LV��!��~�Fų�H��\�����VA�� )�m�b�rP�M������c��0h<?�;�"Zxe��~x^�
�^�hI<��C�G��>��ft���WJ����kI�]�6;:3�
J���BK��f~���WF��ܶqX.o�Zi'Mh�^��Mk�p�`�amO�(@�z�[��Q�_t�fG/�#h�ܞ.��0�]\�Jf����U�֛Qx�cS�E�o&���_\d!%���k`w�����"Z#��a���N%��|��8���q���W̼�7����Cuda���թ�2���C9n|��}����_:e��T�������)�~�/I�	?9�����e�6�;��U_�m�hv�ؼ�r%�����2�挦qh �J�j��j�m�#�"yBܴS��;�^6���t�͎@���j�|Qv�����D���H~�}�1����K���>O�ԭ7$�����4&��dU�"��d��C��k3Bi'��F�&"���Xm	?:�ۺ�(lx,$����<�T+E%�" r���ll�5]�3 g�T�j�a!W��_�ޛ��M:�̦���c
��1P+�n��Qb�_1�7���8����觬0��J�	�h0�CB�Az+֬h����J}��Ql�Dw��#��f� ���
��s���MR��Q�s�j������Q���Ƙ+�(g7N�����D��J"[]k3��i(Y��$�6W0ou��U C�x�-�uf�"��[]���!VZY:�vn�W����x��86����}l��i�+�s����Lzu�!���nnɺ�|�;|��m�Lô����]�zǣ�'��_`���%[hL!�/l��"��H��q�Un��L�R@���~G�8�h����|W�@��]'�T�)P����dbո��};� aƽ�Te��NE[�l�J�.F�&���vB��z��Ũۂh���+�01����+�V�G����DW�M�m;�cL���r_�oǀ�E�� ��H�0���0Hۂ��D�\X��:aN�-10E��g�\�!��{a�Q��P�@t2i89H�^���4����b4��*����5F�	���fŴ�����	�֥[ٜj�w�~y���6\�m�K!c�OM"�oc9��e���GI���� :r�2��h��}x�ƒU����^7xb����:$9?�
��CXta����Hհ�Y�[4х!n�n��UB<3�z�{�˞v��i�^�X,��)^����1T�n���RA�$0���M�҄C~O��e5�������l���J0:��Ox%9py�\�4��c��X^`�tc��J�_�v2�;!W����{�F~ʱk'�q%�U�G �G3�:��s�v��(��m'�:A��¤����(Y����WvU��y#W�]74y���9�n�<B�^�6�g�́�Z�;���6�2�y���մ�Q5�9����p�:_l�=\����$�$PZ����]�{!G����`��S* 	+"W�7�E��EI{�3�ns,�^��//��+�p�q�#��5"ސ�Jϻٸ�ƸB~�
@X
I�.�k�dG�yyU�'�j��(6�)�e��g^��/���ߔfJ ����/|o�ך�(�����o'.$��A1lGFk��LF,�Og?���:���m�����^���ik�X���������r�*�۪E�}�c�����~FR�(�@��o�����ˆ�7&�Q'��O�י+�Kw���,��
�ža3I��A�p�n �W���Ag>tT:b�1���&@1'�E+�g� 3,���6t�J�(s�YF(� � Öfp�,���D}��`�5�g����;��:�X�.��I�����7vz��g1�x2�����AT��9ae�97��b��A~�N^ �����·$��/)��D5�G�a4���b�*/*�+��H[��Ji���?�M3���b��TO�;G���%u�+�Z��b�>5%Z���~��ǲ���NM�X�Q���b�Vm�\�CȖׂ��˔X5�J��hzE�n����<e��Q�9!���p�~z��h��<��V�7�����>�T{����'�AVy�%���[yn��4�>5QFt��%qԏiqZX).0��τ˭BeC�K
��A�g[C&5D��=�IK;�z�����J/b5��ǎ ������U����զ䕒�Ԙ]�k5�h��h^�Yk'ò6?���K7�U�k�"�C��w�V_�1W�����>)�a̭wB�}9��@�,[�%4t��M�����'�9޶�秦�P��� ��2���#N.K~rE2�W�_e�hJhK	z��e�;y��ߤ������HיJw�������R˳Mi	����"H����1�ϴ��E��.�pA�a����Td���3��O�.[%d�2d��A,�7�4�!�����n�s�JI�G��Sd2#�M�$�A����u���:,�.ј�G8煇�߆^��;���2#^cނ���oW5����5����ĝ����
�r���Ayޠ覑N�wQd�Κ6��e�.�p����q��}гCֿ���f{t6�d�u�9a���i��3�+���~HJ�0�i�<�~bAe�� �C�{���Q�|i�����Ʌ��!-�SnrDňt0�MZ�H`���jJ_�GvB��޴��Ѯ<e�2����1�v�ͩ�*�)��)xbp�q��mN�yS����.��}NX�̟�9�F+�\?<�=�[dǝ5�v^�(���T�,���A6���⋸9�<n����G�`b����9��C�~K�sw�<a^���P���x�]�R�(��P�>L����J�#��c�i�|���c�kت�����~~Vd�l2�nP�:ɡ�_��؇΅:D{g�k���@._����[�)�gk=�� �.Y�{6�TL���ju��3Xϻ٧��U@��C8�?:���e���]���E�3�9�s.Hiɐ%Xx�+L i���c�"�|�ϡU�?.�{��)�����B~[�i���,�����_�%t�KP�Af{\��.��bO1�1�Z�و
�Q��:!9�������?(^�/U"�܂z>��ä�
$/
B\��{	��%}�p�(:���O惧3$~�u�v�n�d���x�&���ÿl�Z$$?G�����Ћ
��z?sLU�Kb4� ���HYV,��2�%�)'d��FJ��@"��g��+Cꛞ�N4O������wB`��+��=Z����<�酤�����V��YnT�W�R5/�n�W�gZ.7q�My8ơp�����k�@}Rw�-^��/�ǩJ<͑�����U�Y�v�����QR����B�z����j��A���"WU
��(���c��(^Id��Z���x
L�|��L|��c:3���;X����NU�=�=x���F��N�h������h��� ��i{6��a��d�}ﳯG�s��Et)���W; �)�P!&�V&�mvLx�Ӕ"���F&�<��Yۉ)a�w�M�'*�>4��>�� $�\��.�`e�'��Rͨ�
�{�l�泥�J�z+p��o�o��:���\<�����1`K�:���e����9�6�l9_�w��-�z��HYcn��O�)22g�ko���(`�_�ϴ��ً��w>c�#�?tͨ	�MW�6��*���5�A��u��a���!hC�H:,�'���/����+]PҀ�T+KUx+'X�ߚ�|6E��r�'��2��AfA�E�Q~3[�l[zt4�˭l�sa`�����V����;R@s�������6N�����jb���Ϗ���X�ٸğ~�#�A�:���/��ȩ��s�b�ͺ/���$_�x�T$�Ѻ=�'��C�
�Ȓ�� ~,T��	ZRǕ��ub���?��/(��|X_� ����Ͳ�U�׊!Oʚ=��&4�`�d���ӑ��:Ge��>8��[tͿ���W��X_��[�eydV*p`R匔�`�D����Q�vU>�rw�|s�sFyFa�s�x���z�G�2�bˉr)D�0ף����S+�M��Z�6�M9�v����5�i͸
_mv��Y^Mv�x�Q�{({w�<!$��Ӊ�Ov�v0aYv`�|�@����*��i���rr��Wjh��$����rkmю�G�VJFq���I=�G�T5�6���Fl�>Ppō�z(��w�K����zy���
Wo������f-��ۃE�y;'�=���Ji���6-"R��<4Q��G:wD�~�� 3���.�Fo).a���� ��HJ��#l��	����R���DS��G�g�����_�'��E�8���4�H��o�� ��`d�bc��;�L4� 7V���1�甕��x�uQ�&A�G��oy4����R�@s��|/�ң9��|�w�����վ�	��&��+��H��ʳKq�wq�@�Nw~���k x3h���f�	F�Iy��}�).1Fm��5]"��<dQT��{�`��X1#��*\�f�M1|�q������i���`4���ݕ�-���c���J��͋�4���	��	/\^�б��k[$;Kw��߸w�O���hb�xT�S
�y��!(�!��K@�t�|�o&�:�����t�?�8�����-��Έs�J��R�3(d��&����p<�C��p�z�z�U��gP��9�'�S�^�����L�{;�\�_F�$S$�Of��q��6��+������x6������d��4��0�v�����8��,�A�4H�|�=�]�̢�T��'rM���8z���=G����,K���(o���n��nV;�K��kZBB�j:��/�Y��%A��_��>��*����k��*4�_!�b�Y����yf�9w�b��O��[�(6�*�+�gk��2�������;2/f��e�`�,OD�fD#K�qR����T���ۅ�ZP]�,�����u�d\�sT��|�����g�у�x�k� ��3x
f@�	׹-��"������#�`>��b�A�v��w�@
��3k�6����ڬ�q*��N�i�`���FHx�{2��� �,��w�`뀡�.��w�S=��:�����n���j��ďx/l��f1ۿ/�Yh��a8rH1���O� ���Or�s����jO������̡Bj7P�ȷ�0����&����DfvЙ<ث˷��k�.^�I$,ٟN����ӄ�sE����PY*e!�1����r)*�:�E����b��5_�u��t�]�lr�wH£+�����Ղ}0���VOA���k��W����`�u��ݶ��{vp�v�K�,b����K�+z�4��a�a0���+I�\8���I==�����U�]+~��OaR�^�\������f�rf������ä;�N�L�׉���y|�(��\��"�۶:��A*��Ƨ�[�5��7��znM	�:�e1�"�拎ة�!�'f.ʒ��,18Z�)2On=+�S�b���j!��q�&I�;!�ٽ��v$(�9��T����irč|�����h8kJa��9@S�gYB���2t�b8_�u�X�x�`�_�L���F,oj�R���1р����D.h��vьL@2�6w'G�,����W:��怊糱rC��?R<����m����Â1A]D�n{�z�v��K70�4i��%�oeD]�2�ev��}��B��@�.V@(l��A��i�h4\�K߹A��wO�uM�6�w�_s��z{���vO�5�Y6���	�.��$~�2-CK�}2O�ޕ�m�Q�i�p��=�(/��kf��+Ђ
�.�(CamyJ�����Uo��"�Q���Uu����� R�����/tAzJ�.�n-��ه[�]�ͽ$�L�`�ip����2"���n�Gk���d�B*�_�}��15|a�~4wX�3��fwj{���,���+X�c�|��DYZyU�R�u��Z'9�N�,���7U��h��D�4����iw���@�bJ�х8�?��y� �:Y����v��3th�)�c��3[�2G�S� ;��<L���"yQ��y��\�I�7NYt��i��?������c�My�a���9�F�[H���+��9	����JѬ.Rt�1%���S�G�`�K�01*aX?T��1(��Dõ�д�y��
V�����c�U]��?c,7���e1O�0�.n�#�?-v/7�I?�T'�e9<���f?�[R�:�����-m�3�E�+��3Ŝ�m��a�=&��� A��O�J���~x�-龋�C����j�GϘNT����Ms�-�΋[DV�i\���h^6̼�Gj-�� �j��]oޗ��d-l��t�Q��.r_�P�p���������G�^�g,+�a	{m4aQr����/�����y��ϕ#�|�oX9���o�w��H<���Ox��o�(iJ�L'r�q�%H@�y�sU�EF	U�vb����6�Q�(�����'�����Ө��@\ҹ�����kq��I3|�c�ų�?U����>iD ��Ю#樲9�SbJ.�wwW{Q�Ra�#z��R���ֻ���������ɟT���˕E���A`�IEKȻz���3�{�`6I�
��z�8h���'��  �6X���>Y��ޕe��@!���{z�Às��W���=��^��4�G(c��ݛ&o3�=P!� ����i�6��#	*kn�]�l�>�;�	Ɂ�0;��j�`�k�O$^^����2&"��3*��nz7���V��R��+.���~~�R:��Jh�j��&��9�ɉ���A؄���Z�+�2���V�T��2h��ѲM�zP��P�b?��G�?����|Ǚ��E`�ݽ+���F��:���i5��O� ''W��Զ�����~$��8�"�y.�Fy~���A?�;�5�|5�
Z]���L�x��Z�X��*Vz'#O0���׸a���X̉��!�v�(�\Z��G�Ҁ뾣�w֙�Խ��Z�� %�|yq����\�.�r��D��UP�pe�o���>��6�fրN@#
�rB����K!�ݯ��l�����)k`��Ѱ2���R������>^ͯ�7[-9��,#��Q��� .��P��I;�6���S;�zF��AĀ,s���;�TB125=����I�js�����7{� �bd�\�Ws	=;s���=�پ�0aj����f/~D�ޚ��0.�͟oKAȞ� ��{�!��V7	�B���5�H�R���p-���b��s��z���D�9����v�w�z�&R��r���B������P�$k:㦨E*z�J^_�H���R����*5��� ����^�d�A�k6���E;���U�R�;�1�������|(���޴����1R������O�]�@����e�g��,;|�}U���dG���1;U����� ���ϕ*�]4�9泷�'���o���d�$6*�e��Dbv�5���;5���A��������q����]�t�0��| �L&�"��~C�/����6��[�cl"��n�zM!!��ӽѠ��"R�	�Y!�������B��hOfra��l���W��W
f��vÔn��5Ht�e��^����o�A' �J�E�)�L�b�B#�E�.)(�f���Y}2ʹl�!P�
����0|��-���_��ރb��d��q5|��3�_M�m��E���� Hi����e���Ƣ�L�X8��z�ul�Y׎�O�!���)�Z7�sس%&Z�G�,�?,�}g��Q�(D��\77�c�e�@���^�i�u1委G�O�!7h��ÑZ�e�_92q����� ����Fp��1g�so����ʝ��C�Q�62�ew���/��)W���7��}(����&�˯B�5�\]��z4��k�7�>V��r���$<��@�3nֵȪW����T���զAOI��2R��hϿ�ri��gSB��>�Mr��N/ӷ@+ΰ�ZC5�O0��l��J�����0�i\��d����QP�>�ku��3�֟mQ����/�SpZ��Ld���l���-X@�0�ta(�6dk��U�U�04 ����}��`�Yw��<�3��Ƒ#��$�S����`치ޞ��`=E�lݶI��oh������ڲ��mz��V.s@�џ��b�f�V�wS��!�'��/�S��C���^�#�cف�S�T�+��w�B�qm�2{�2�x:�g,���0m�G�KS��$y��ĳ�|(W�#��2j��~�z�_(���*Acyׄ������R�#̍���an|e5'�#F�b�TF�|=|Cr,`G��ҏ�b��U�/��I��K D�ѝ��C�\����4�nV�j���IlP5�Sm#9�G)�D�嚞�ؖb%n���Yxp,�F�m�&������C�:��*��\���ǋ����o�N&���@��G��r�{�b
`W1VӅ�~�aO�y��(=U�YDP�Rr� 5F'��OhY-h��Ⱦ�Er���	���l�aK���_��.��6!����+�1Z9�,!F�$���ov�nCV/�]�����705X:
2����7;�Hoj`����f�G1*�ȟ,.gO��S��fE ���,��jWz%�c�N�	��f���3�����#���O���P;&���JA�1l�֙r�|t_onQ��V��:Cm�&�lU,�f���n�)����[�΃/��Ɋ�µp�*��2�7�2��c{
����DT)�-k�;�@��u9$8�l�)�RW�S���ĳ	�qa`�C���퐨<��3���	*PƖ��g�VE�E��r	�6�U��ז~���d<��	-��m�Q�N��1NHz�?4p��g�p��-)��DV�*Z�
3�Sv���c�����;����2�I���y��c%R[��P钛_y�G���1�BS=�1� ���<�Tz�qN�X5�6�&��y�ݨ�{A!W]���x����Vf�;k2���Fc���\�	�� ��p��P�>�������5��½%��	�ˣ~-3tRZ�v�>M,�j
��X5H��zC��ac�}�Pg8 �p��N���CL�+� �hS"ߡ�;G(B����C�8,���;��8��T�$lA-#cE-Zղ�&�i��X$i�xϤ��k�1�&&5� ����AB��czU���b�|���"�W�m��
C��8}�"�n��U�&A֚Em�y��8jbtR�	pK��T@3�V��?}�����k1�1W���.�|e��O�4��3�	gp�D���t@���5�ʄж������R��5Z�����Ʀ����Ǝ���F�2�SiQm��>��%���(y��؋.In�|����M%DMs�Y���e�_��<=|�Ï�㸤~1���631�Wʫ���.�m�s��ǵ_{\�"���ȁ	�!9�7H��|���-�J�����,�����3j69lY~�<�ڍ셤��)���?=v��P��.B��m����AA���J�9%5s���qu�&M����<��X&�|}�d|e�@����J�.
5I���W ��R�`��#�nk6c� p��V���0x��j�n���u7s7�0��>�'���
�;�,؛��	���%��I:��B3~��ʽ��f|T	�p!p���C5��KQv�bG��
I;��gX�fp"�s8����z�,��(-!�&i�7;z���K�7Q���3��\�0��3��
�i�5ɕ 1L�pZ���9��8���謻��--��&E�`!�b�5�+t�s�ڸ�r�s�s,����;,�� /�ŀT�jL�f����{ �����/[���W�ă�F8I�Of�<$VJ�20��B��HUOLT+ZJg��F����!�Y��N6��&�B�.�e���!��ZxL b����8�Czil��Q��D�#)�30)�^ó����
Yy����6�x)u��&͚�ҋ���.k(�`��Z������j	��o���d�=�����yD�2t�x�@�iЮ��9p{x���_6�r��6u۲��t�M��.>`�.��t�ҡ)
$������9�A3��">` -��%�����!����/��1�d�g��%��c�eg>yVtʺ�=�#0���}��x�V�e)�DK�&h�G��ol-v�*�ϝ.%E�'�Mre��P|���"�f�|�2�gq
K�z�FF=��S�7�q/�%�5�\�m�@�IRbrj�ב@{� ��bN�7�q��
��K5�����S�����-A�F2� lD��l� �˓��C�c��U�H]���@9�,�W�[�Q�C^o0��<�E��_�^}&0�8��!NJ�7����;�j<?��!܄��KC����.���ָ����~��+�T��+GP� >��+�Ac�꠿Ĝv��9l�=��k�UPkv��ȌǍ�N���"v��a�`_ܕB�����繜yT.C�>�=�=���^�|�.a��$P�72�� ʿr�z����$̅GX�#Q�^�_G(�C�է%���_T�����}��A� �������*=">g��lzG�_�i���jy��eBӹ+�?�[�ɪ2xOI������L-wU���A���8����A��q+��PA�2�޿�3;��o<{��5�L花n�y�귞�%��2z���*_�
�[�Z�Rֹj̠��'�,�/qQ\g�5T]�ۋ8�)3B���0@�q��-[��S�=�hϚ ���0
Cr ˇ}������>iqP���Q_N}�� :0'���Էl����Z�j�XAFu�VrcL�o5F�)������2n��A��Y�P�e��|��Ž���R�y�aP\�D���K�Ss_�0����ck�å�u�8����U,up,D(��3eKX���P�_o��r)�v/����
FE�wqډFW9� XC�?�"x�g�����A����rS�� ¢Z�����ǁO��O󚃚�wqSv�z/H�a\�7|�7�bd�0�p���5b�r܂�^�K�)nRق�:��̂���lԐ���$v������2�F��y_��s@��.��t�??���=&s��Ҏ�-3��K=�on;j�e|zt'e^0��/�󀳹��#��ofF�$��6��+��;2���10
+wbRz{N,ڈb�B1���e �ҎՍ�����֭cȮ��@\�]}�흛X@x\)q�g\'f���%�I����7I7M�n�L��~�Yp���Mi������kyq�آ�nƥJ͇J�N����o�|\ٷ�ލX��$8M�e��>P"H(vg�	�d�LZ��j�����n�H������!x�-����|]���5��3_��H�.��\[��kiP����_)Mؔi�4f:�
v��X�D"��b2�ҜqӨ�x�^��������r�'�A��� �����F�/'t7�D�cR|��-�]�mq3xs���"��eV�_�߀��~��� ����������������Y$T��8'�p��X�.���ͮ�I�n����bq�����EC@=#T5nfhÕA�Y�z{�b�=ԕ'�K3�t������ h"�1:�`�_��$,��c@/�[�a�r�t�)~����!l_C�g��<�ҩ�w�E+3^��[̈́�y���sj'~�':4`����W�Qj�/4�0�x�t�ZqOdw�<�+�!M��ܔ_\D3���,%E2
�*�M6v������y�G��W&�X/2�
��/�Ӛ�8E�Q��?�e8cײ{k�@H���=8��3"+���Iـx��QG����/ဣ�]h��<�dfY+S8�-��Mh#�?5�a����T	q,���ѫ��N��14X!Ϟo�Al�Ѹ^�'��^��El|�0o'��y�Rθ9G�YI�!�L�)B��{!���j<]��H�0w�/�ǽ偟W��_�c!=����g�pK%EJ+|��BN*��i-/t&�/��vpC�4��^c�m8<9(�Y��t�x�74����� m.��.����*��7����ν���l0M�!8��)zl##s��>Q�ʭ�P�G{��Ys��KY�^e�R�o�
\�	H|�e�E��)�D��t7]�7}4k�^�C�X^`w�������_y ��L,у+b��G$�ҫ�]$
��>ĕ�j;0�D�#bs��zW�n���K���� �	?1���%Mߙ�f�ār��KE��`��j�^�a��Bڰ��u���xx�D/���뺥ٟ���o�4��[?;Ҷ�$A���:�+���4�ʴ#����Ǽ�P7&�K��X#	� _|�?T�_��"H�P��t��P�⊱t�����Ӂ,A��3#1X��8��ſ�a�i'�I��U�@s��}�IY��Oo�;Y���>W27�~ͽ�+^@2iB	Ġ�(sU�O���?����n��6�j0C���H'.RH&���|/z]�q�ܶ1�h<\o�{����xNK��L�c�QY
�x��h*S�e���O}�9�ܤ��� �J�l��ɍ�+���|�)w1��&�R��� D��A�w ,�b�[Pk:�J-6�Sc�{�('g��pC��A-��IfW�,ޚ��~�U�.�[�[|�i7�&Na�?�����J��~�qG���b����ӾVJ�2)�3~��S2�
��ɝ�!aϽ�#��~�Í��W8IU���,G��H�^��28�$ܡCHAH]���h�oE�fF�����s�Q.��}�r���iIB��&���(�Y���K_�'�e%��b�N��#/_B�����P���T��L���k	O��py�4�c.Ӵ�Pv�܈kLn2SRP�����4}��[C	�(Zp�&W��	}�Bm�b6'=E[Tu��i�x)^�4��Fx���'��:��+�;'��7il)�&kY�v
��f�ieV��!�uW�?V8������.B�19Evb�E���Go�X�dZ�,����L�
r:����\<� E|?��"`�Ů;�aP%�h�y!�+([^���q􏘔�c9�G�"��y�'��"�piE/w���7�1R��( 4����&sR���Ŭ�MB�23���A���฻@^�a�vԐpdo��Q�`eJͭ��9L�6F�i��+ҕ^b����*�ՃWTUS����u��y���X�I��[��n�7�]t}M?��ѐOթ��O����錠C��d�Ğ2�FL��L��FZE�K�bx�G������[�����������,L���r��D�`ET ��&��|�$RɓѾc�*1b��AYg'��]D�k�x�)�������l5&_�Z� �ߟ��2%��.�vJz;]��C��~�Y-��c�00/��a7H�k�z��W͹�w�3���:�K�u�:d����]�.��e��|����#����)'}TC�R����	��Q�%������q'���";`o���M~���[��:,�Y>� w�M<ԣ<���_>��\�BtI�38V�q�4�`Vm�2DX
 ��pB�ϱd�<�cur%#��X8��5/���@�k����)��g�e�!j�|D�����AQNw��7����ߚ�`��˭���a�[�#��W;�k�2z�:�F�� �%&R��� ���Ƞ"�zq�%
�k�1��l�{ h�eЋF�k\��B�iqR2cH���O�'�;(�.�-o�S��S��I�J�> ������i,�p��MƲyï]O����T�'}��@�z(Wve��c����)�RC���5<Ȃ��M�s4�a2���?���%��pW��.����
]�����+�e��9ٙb0���	r&�-�F�?��7��*��&�i���8܂g-K0�(c�Ue`r1�b�J��}�;��@6�`���"����f�q���x�u%����z��o����'��`$ۣ����BB��x���dV#2�a\g�u @���"�=�jۑ��s�/���@n	N��dl��p�~3���~�L:�<:�i�:�b�(���	�:��X�^^���O��TB���S�*�q���M��Y0��A4�1i����j��b&_��ڐW=�fY��y�פ'�aN��MԷ3D��+�ʶl��!�@�Eq�Pl����z�M�j�O���V�D�\��2��0����,� Y�;���E���}q@y�u����~�/k�Bt�3����P��!+Z0�EQ�x8g���"��G��ަ�ְp9��
���K?c�~xnH0�j ���6�*���R�m�91z�{�6/9�6>w���F�#Ki`T-9��eHo/^V��'\@I�������A��y<ٹ`��LT����Q:�-��;������w<����LN� VbC2��)�u3[���ϲ
{k��|3�?D��������HN����<�P}H�6�v ��_?AG���:V��2U}�I���%���_	�OcL�Va)��FC��>�4�Ʋ �[��*:Q��{�Г�OC�-�簳n����z�ҩ1?QX��,�pg�pH��`�?�;4��I@���ej�(��2�U� ��V�Z�|��d���6���8ȇ�C�'��z��%B.��/��S����h=ֶ���Ϊ��F] ���s���� һ���-#ePJ�)��X0g\F��Ctd�&��6&P��C��h�SĭAX��֒y��0�vO�Ш�J�����:qӿ $��!%�!�Ar$T���3^B6�Z�4�5ܔ#2v�T��4���A=���+LE���<���<+�V���'f��9.�[���v��sf{�D[��X:�O�&P"f"��tH��:�74Z#ES������RA�F��>#$M, ��vG�n�E��6u�'v�y�ύ�db/���F�!���G�ayy6��?�t��C���k�"�<z��"��gy]���sW���ZPL��Ҝ��^=_iUw���9���0m|�x>�y�;�=4����e�g�P0����EQ1��`�\��|�n�A���� ��"ڞ���� /8��t��0����g�r���k,3�L�XI�_���L%�<f�~���66:���,�2g���'��bn��R� 9�s�j��y�{���gD��&���p�ϛ�������xr55�,�(��L�^��s"
uPq[����z�ۨ�'���+�&��}c(Q����;Ifl)S�MZɥZQ���PV���r'��o�9�.�!&��d��)��������#9�y�����n��~I݌\\i�C7�z8��%�[����<�ޓl��F�~��M��}sN+�o��^��-�b'���o2�sì�Us;��#5ÉO��r|�=��@�q�/k���V;@�*[����9�I��^�%V*Vf8�/^U�C�.2����������2N���cN���Ŭ��ae�b�I-VL('��n�=ƮW��B�����=���G�����<�0��^�mf��V�c���sg��ȃل,afkoТ�����^9q����tA�eE���jA�!V	��Nv�z�nz9��({�:ke@�f��~��om �{t%<D� �mW/���c�陙��p�ﹰ��f���U��t��_�|=6`w%ۖ��@������g$�^����ڸ��Z�ڀ�u@���ܿV�cM��V���� ÷�3"�D�R'
Q߂37	.
�-�'"O�v�Q�v��B4�x��<8���Y�.P͕(C˩]�����IZ�e�Q��Y!v7�P�]�Uf�t:�Ѕ�i'��?RPfJ�!�?��Q�H��ME��K�h8�Lտ^�eW��Á�_�{����<ҡ q�|�b�W���"�pO�ܻ}ô;FC�粏���_���ε����U��^���yω��K1�໑�˥�@4�(����m�Q�#S�O�R����2�<m��H'�L�+H�?���u|���d����̇ch�{�Z�%��$�V���X{����X��vƍ+�8>K����?�Pk�"�y���''�,C�/�;YU'b`�ęrt�E�����C�H%����Pb����\�d9v�M"�Iu*�w��8�I2�!e�S���i�S7n��l��
�����rC�ؖ�� _���.�ZA(/3��u�avdͭ�h���8��ѭ���y?[R�ڿ�S��Z>��)7w�sȠ�b�#�]6,�/͐��w�^�r�=1�������bհ����� y���k�s�Y\���9g(�˫�9�q�0O���)�G����w�����xG�\�m'ej�T��v&����V�C�l�G�h�eE\o�����'uE��Z:_=���WE�2�}w�9�Ү��&��������1�)v&U��?,�d�AqS���z�ޢRv7G�ku] ���%|��Ĥ3���=����0I�I�M��g,x���,���63�A+/��׈�z��S�q4�wm�����X¯��ז���_�o]������
�hd��?��G5�m\��,@G�=��o�	8�^���/]p1����ӽ�u�E{�[�=y?�
y+�xfhmF=���`�_�W;iͱ(Z�Q�d���P���r��I�.�.v]�� ��i�V,���tQ�W�����)���}E�c,ynRS��B��y# 0֤z�����������ߔ�N�X@�����1yJG��p�}o5u_9:����ǮѪzi�Viv/j�����z���mΛ�v���޶��ܹ�sc���W�9R��m^CɃ�@Ŋ�1�y��Y�\be�k��*�J�6w�}�mB�HNM�Ы�,��W�e���y���RÖ�d�:�;V���`������;�@�����h,��º��mY��k�W����QY,�՚�y��8Yd�<�#�8,��/�����ld��V/���L*�̼�<��K�v뻷ΚZ��;x2�|v� A�{�.��h�տ�H�K��[<��fY���m�KHw<��	k?�B�4�x�J#+��3�ܸP+���I}e�agD��b]0��x�l�V$rK��ɼ?��k����c^��T��J�H��e�b���ڜ��-m
�cm�s`�ʊ�����w:졝�HaRm��ܢ(�
�!e�t�Q�(�!^���j�~j��5�k{s~i��xB�w�F��J�R���F;�'��������6f��K��r���)fjYz�O���tF4["�q�e�\U�-��9V|�!&C���E���H,�s��s�s#,.%ͪ�M�>A���j�%��*�x]��*axt�;Dm�ǌ�#Ge�NR�=s����'�^��d������:���� �Q'm�oz�Rk�q+S3֌����ǀ��:Ek	cS3#&=_��/}�ѥ�*��j��/-t�J�+fN���D^>���x%�B�#��Tïw��%�D�ti	�0���cd��
c���v���H �w�s�f#Pi���o�k�6v�'Ѩ	��N��i�XA+ZN�"�-��s���ǂ�RmZ@C��u���yqt I��L�0oBeeim�@Gs�������Z8F���U6Ë�UK �I@�2ⷘS��I"�Ɲ��G�\� �z�������Ȁ��35�A��A�?M��]΃I��d60�s��;�̝ )Ʀ��]"�/�����|V�~����T�(�i�u+��K�2pe��4N{	]�=eo�����k�Ҷ�[������~^�9��T�?j�'���� �iȰ���+���wT�Kr�S2M���?�@�������c��>��%:���C7�Fׄ�4�*'�.7��|�JT���|��/h���8߫f{K�[v왍y�z��d���'���������!�i�1�\�?�'W�x�5�θ�9��_@	�@4�_�+�� 8iz��Ս�Z�9�bwV�Ej��v�H;0^P�o~�å
"��D��G��6��������2$	$䬎��{N��џ�����̩�;k��/E\�j����G:�y�'��j�*�!���������v�D�L�60�G#�� ��DlE�:�J��2W�d�����\�ϒe0�42 �F�N��!FcS�9�?D2uy��vVlx�T%>��["��%��)I�vFk5�ȉ�]�%m��2n��k�� s�Q��v�$�G�wdvt�]A��h�_�����F�'�u.�Cm�l/��!����Ƨ6�K�Pd��7�o!��Ф'>�ZIo���^&<�~L��P��V�/ܶ�a����0C��HU�g��?]h
�f'�1t��-д�4�n��Y�����<԰������b�^�a� �:/x��K&/V=�ڗ\[ZM)�x��m��:U��v[Eb|�2���}��()�~ph~eW����`�M��c�uX��^�$�n!0��9�������/SrM�#��/pn�ے#�_�q�+�M7P�\`~��1�7v���hDr���ܦK_SKD����;z��y;��H۵*�(\{x24B߈�6T��"x���U�$�������,t���>�RB��cL�Z� ����ԋ�(��ʧe��,F�y��%�Z*|�Ҭ9OJD�5P{;qhQ=P��ͷ��-�z�m�Y��C�	�b�f��G�?���C��?��75�6��"~[��V���J"u�����,krn�v*���o"�N� {O�z�D����n��o���DQ%s6<�L��7��A�m�*��V����[=c�����̻�Z��6M�?[54�x�{
ʇ(cG�/�)���� -Fa�o2ݳ��I�	^�_�Bе�Z�Ό���n�Q����t��FI��_6�
Ι��?l-^)�
0��5!�rj8{��g�;Wc��
@�je+	f7�i2��H=�VP<��k�D�v�Jʏ�,W#E=�X��g@r�Ө�9�1Y�{t&�oٞ�NX<�a�D>��?�_7_�C�L���������)۔%HRq�0�뿿x�6T*e�ze"�r��k�.G���H����2ݱ��;"��Z���[�`|�C��&@��{���&	 �2P��aiE��+�9�X?�>�i_��[�:�ҙ\�	'�c�* �ޏ���CF5�=�EQ�G��_Xl�TZ�����*Y|R�� �M������k �W��.Bx��0ҔU_�b 9���_��;=�S"ʃ�*cq��`�F2�i�Q��,`��'������t&���?�q���.�:�t�a�� �>��3�p	�	#Τ����^���tOΦ��'m�h�A���r�$�E���ͦiK��z�1Q3N�:�,*F1g:����"o��=J�v���2*T��i%��%�:0dT���W�A?��e$��M0В!Gj�鷰�'(���'O�8͛4����0�Q������R����4H�X.�g��w�9�Ugp�Q���=��x>lw��*g�W�����}�A7b�$�w"{�ہs~MX9j�u�L��含�xT���:����i��4�Q�@sN{�5�2Q��!��R��?��V�,�ꇜZ3�u��X�h}��M���\����G|�x���.��C�J7J�h��"wv�jTꖺF����ߎײ\�z�el���oa��v��=���,�s��$,P����k%�6EQ��3\4�4�qK_��N�x�; ���N�-�c�?��<(s"$����<�D�[���{<e�@(������H�5��6T��R���JR��燭�gP�ٕ��?���Ѩp����}.p^�,��	����f�@�	dv���Ri��O~���-0��zU�X�R�i�O(��6�бQSa1߲ϕ�%��{N"=�1MI�Sf0Y���ܟ��\ڑp���8�s���hw��oٹ"c��4[�3�wU��K�N��r�a���?Fʏ܂%.�l��=�!���s�RK�E��)B*��	�����T��*#
|`ɱL���v8Y��c����Z��QP��8/A��I���͊Q��v��ϭ4������C�)XA$�jz���$�#���L�^1"�G��)�	�jx+=/!(+�}��f� ��<2�t�,I��/��S�2�\����jp]8�(�!φDBhd��Y�S�%\lt�{+�x>�����>7������,��_,Q3k]u�R�>���@�@�"�)i76����ڥ?4���X�j:�m?����m�����Nui-�,�b����3f����_�o��]@]�H+�7��L.��-w�7�S/�b�����i.�䋶�Ӹ�aZSŲ��N�Of�]͓J���j��p��DŚ`�mĩ��Q�����.�6����!����*%��a��׭��x��߻ƀ���sb㱙��Ѧ�VC�#����7<�a*��!��=-]�[�E�M��O�jG uEi7��iw+G��N|��&k:���
"��u#��-
����&��k�c�������%H�_̢k9`��D�'G��,���x$����+Wq �BBe�`���� ���$sh 1#�ǣ���&�L��$��Ylvl<u>S�0I�$�Y=�V���s�+M�+J���oG���+Th�Az��'�H�����7^�}�qa�>Α&��
�&�����u�E�	�-�eGI�SkXF�jȖV��%���y[�}�Ʉ0���m1��h��~��$e<l't���~UU f/SM����e�"*Q>�K����T#4U�F�d怎ޘ�69y#�-'H���k�N<�x�4����t���@������8G�痸ϩ�8Еp��՟&ԍP�������v��_�)1Iq?]��$��l��<�J� �q}��'Kj��%��m�\3��9��Y��s)��mm����m:��_"�sZ�{���l�<��B�R�K�A��"�[B�kQ���rl�:n��	^� Y�O������c�X��ڿ�{�S�����f��xz�N��b�Un5/�x3{��\�q�?[&�>��寍��$t8���X��&�S�����
�����'��h!q�6b�٘ZL�~����և�ҪU�n���ܲYә�E2qg�U_2���(��32L�SVqG��L��*h�N�O|<,"�����4f/eь�������&!�o��%�{�/dlG��$�n����;[��3����X
Io��;�����V}ū{S�yߣ��<%�]����1���R��I���U���>7w=��h_�4�&HH�Ja�?��8�g腖6m��(ǚ8��g�~I����M��I�����_�� ����9�!��5jP�B�TXs\9�|��^毴�Ic�@k}���6��+؈˷��ø������k\�2^�W�F|���c�	����{�lC�Y�Zʬl]_܎�V@��Wv�@)�� `x\ʕo��Ԍ�,��X��1�>�O%���d���n>m����t��yw����gu��,3�oo{g4�*����W���H���(z���w^c㦵a�q�B^��W�3E�~(y��ZV�0
ִL��x|{[Cm�L8h'��I�-Z�;Q}����Y��0@?��ԮϚk����8��j�w�י�;nX���-��;,��ƪ���Ֆ #?���}*;6rC��X��j'Y����%�/��~��j)�*�a�"� ��}6a��6֩�F@˃�2��c?$,
���K9�ht5e�"��F"?�ė��}N�fG�.�G1��>&�7+Ia�� �7\Tk(F>�	!��g{(��ztK'8�Ly���Պ��lo'kF:j;��=U�J�h�JdzN�f��QsX}�i,���j�^&�?fK�6�K���ip���iA�M������F�:ȃ�Q뺶ߋЇ�
I�[{߆�s�$����U�T��/�P���fx�˶2m�YRZ�	����l�Ql�T�r�~,�SR(/.s4!�,��0c�N�=�M�N	����1�|,�(w�-�M��x�� D-l�~˪�P���TEL�-�rYL��	��n���y��$���,
�R]���ص�;����o�9]�Ě�8�+��|��
�OV�j�rҦ��-�s!�f��SJ��2�U���i�����2\��3{�ӂnT����v.t�R:���=ޖ]�e�K|b��F�s�;c��m��R9�(8i�D�fbq�:.�j��]l�cq @����{��Qtd�;��d��)�L�-�F��v<1�X���(Ɯ�����dW�%f٫��,�&���Ґ,ר+��v���)��`������Ov"s}*�(|�}ҍXOm�	�J��U�4�cI|��'�T���Y�;�Gj�XY�0uէJlY�3�Y�Zc*FC�}?��HGH�w���MƔw�N�MlH�i.Ȗ��3:	�����������A۹��r7�*���sd]�D�]��/���I�ؔO(��69� �g��O���`�����.T"�l2��I�t+�GN�!�4P������ġݵ]���G�������y�Z��<�*�;��$� #*pO�b�e����f�4���}�-~O��j�[<t�	����1���3�|+�C1|cz�1����P���e����J��+<&e]��=�/��,������^����i-�l���X|H�o�b�'_|%#"<x�20SI��/
��P��N ��i��]�h���}���hHU^&vY�3�ng�,O�� |K��� 臍�@��� �2�`'͏on]�a���mOQdp�S��&��͛L��I$V�c~��%G��6lW1	��ꌎ��du�� -[�}�2 !�2�2�ؔ<���-f[iث��o�@�mwG�~o�}|���T�{܊�,)0	��j���oLg�r��w�*���g5-Q�ѫˀV��Y%��۫�K������`D6��z�yl���o��|�SpP|�o[t��.R�'1�~o-D2l���K�` �?)����'��~��e-^�������+�C
� ��Ld@��=����U����fB��s%��t��<1"�o,��7X��%�;��|�
&��d�e��[��>ҷ�6�0w3�h���I�wn3ݧ� �b�U��4��f:"2����m��e5?T��E���辘V_KH�4�.%�CCq��J�^7knAv�V�N�:�O��Uұ>���ܦ�Q��9"M����l��+�:�̬#�� 19�웑J
�>vGoŒ-i��M��`��&�PI�z���{���?8�y��2��C��h���>��zb붢�AyU�I?3Cv^��� ���W,�8�hO�d2����s�\U@'���ĕ�x��Tz��j+T�2�׾W�[i<i#��`�2�.(1W+Wt�Єݻ�|޶5�R/n��z��v7o��um˯�}b���(u8w� 
Ҍ�j��|a;����VRs���z�뽸����lo6�-�����g�.����#����U�ɞ�z��VRWX
�(%����[�o�y�X��o+A0�s�0����+����������!d�){֛�2�6�|��-'%��>�n��`�P<׌Һ����E� ��{R�(�<���t�	2�~�b�=�"��_]/n�_Yt:�@��]��
ѥߍ�gx�E̎��%)E�Bs�����L	��)�LW/���x��`�3����{vL�\)�Hm	��M:@P���Jٗy�[����1�� ��6|��Ј.w��! �gS�Q k��i�%�Ѵ:ߘ��R�N�T!�É�&-�>�9�y"�����|�FB���J.i��=��b� �i�wfB-Jdp$� /��Y"��� ��m]`#/ɫ0O�S�p�h� '2R�#!K@Z�]۪��cn�,��ݟӗi����y��[�5�ة��_����?���Ƨa��b!0���Ө���C�FцJ	^��{98����Y�H��, ѽ��Y{ �55���c�p���ȍx�����T�񌕍P�nwl���dZ�M�T����4K��j��\�Źr���Z�
���&KZ>q���5C��A�^�s܊Ȋ�NΘ��cYm4�bd�*�S�ԄF�8��g��}~@{���'�}�g	�s؅ �w��(:�
A��˦�����2�I3�W�?�q�~�b���=q3<*V�/��=6�es��r%��X�����F��t�ʠ��*�U��/�� �m�C��ZӘ�^/}:������w ���F�Ӧi$E�g=d��8���JH���
��ĕ��5	�X�}����R�w�H,F'��tn�<���ka���aL�*g���V;���������xH��B��&h3d�;%�^���!��Ta�u�y+<A�`�Ƴ�� 1ʦbgM)�l�':yba�sE�A\�$�`
�~R[)oҏǳ�nq892�>s�)���հl��ݐ���Ay;��`���cbm�n
]wsC�m�L_�Y���f��y���� K~`Y'ޥ},�6��?�6&V�;���J$�/���|�$��ƨ�,�b��ޟl�uӚy�`��t�H:��c�� ���P�+�d���dP}��z���&(	��rS�ڻk0���J�T��2o�>!촙�-�^��1h�j39�9	��p�4�Cɋ�=���=�4�����uM@G$�k��������Uq&�V�!�s��`1UY!ʹ�=>�r�������}�.z�eG���H����e�В�?�lL=)âf>�!?�E�ʹʈ�$��LF˨�����B�5D�Y��4(�2EP��χ]���ˤ;�X��Ē�o,�\v��:��^�����tM�ho<�ȿ�[[��Q��J������¾�YI=I�����!~I]i�8�9��f �ҿ�dͫ)��pu��yjr�.�{S���3�ʯ��1_yد�n���t��f�-M��U�Z���x����Т�I(mW��fϔ�s������$0��#�+E��˧(��I��]���׀1�r���]�~NI~������]k&Of�n��CR,<�-�5����9)%m�F�[ⒹJ��-YY��#���^���Y�&:�j�������K!tȲѱ-�Y�>ip�/#<@�8�j"�	�z���JSW��u20�C��-�_ڔ�׈�=�5�ڒ�czH9U��$-��M�%�u�4q��\�y��4������\����b�qMK�$��3F�ީY�� �����	 6n(��f����)8n��Ӕx����tb;{�����Hx��~��y���|�>l7kf'��M��-�6-��}��!�iM��'>��&����x�cz��7��0L�$�Z�֜�56�p%B��+!�E �Z�"撊���P�$�u��հ��׈Sĸ���s�@qV���&���r3�M+#�t��ӈ蜫���;퉬D�j�m�;��jFYQ�4Ɠ�;2���eݤ�vW�ћ?�[/�o����M�Bp�)�M�	C��C�\6���5P�*eߤå.ැ�-��"���Ⱦ>}5k$ъ�mƙ"��@��g�]�B�z�X���pT�z���_�6B�V���j���K� ���9:c�փ�(LV �;t5��� ���?���К���Z�+�6�ed�x#[\�z)֍��h�N���N��?P*$��#Oʢ�G	��H&c�1]�g�����;gdd��-����b�4c�#�" a{�ԕ��|#g��o��Ђ������S�@#L"���n���g�yK��UGȮ|����"Q:8j��On���S~f�r��)��WG+ݘ(�3�w�{`#-��Ċ��\�=?���_��_8:?�,)���j�)�ڒARu;K�a4E�Vm�M�~�l���0�m���݉&� =�7����?z�#L�t�b9����f�2�3��a�hp��6�d��O l������E�,؋�
��r̶��z��M<����d=��G�d0��!�[~��E@T����1�a���Y)dּ�*��s��u;���]�M����,�n������DG��LBn	���^�tlގ�u�jn��r�x�3�sH����1�;����
W��Oɂ�]�Z�����@�����3���κb'�r]�L�[���A	�$�'G�U�������	����tG�C�"z6���/X�;;S;�ڨ'�;G�K�#$���#�s[ez1m7�^ߋ�y/ǣ�ߣV��p�*��v��9�>0����Q_ɇٗ�1"�M=mbe�j�6U��>�}�#�=(� �FA��1hU<ѐ��h����i�F[��!�>��I�YȤw�#Yg��0�`Sx�<{�@r��b�3�8"�W105��+c~�y�a��v��x��j�wi�F��;�s���[뺴�
�k��ʬ�N�f�#]צ��$]�@��,�m�aq�TT��D�'�s���I�W� ��$I�0*A�w��_)˯W�li��1hj5U%v-!81/�zy����_U�[�f��4+�M��0!�H��t�8�#���邨s�͙P���5���ɸ��4�ρ�8�#P6�v�0\Dh����M2f��F�_5��e��l�\�u��������#G��|Q�s|�p�k���)M�N��FY5`a�D�6�|���teK�hV߇P����trh��7��k��M+8�Q<��rŰ��m�/liޝ�$_>5�+����TV�2	�u�.Q�V�߁R/82a���,��7�.�2�wa*lvU2@18���@ {�dH|���g�P= ڨL?;ȳ�,Et��Q��	����x%�8~�&[=��8����*g��1OF/c�/�n9��V-i�nuP�.a�}:� ���F��z�J������Y�Y���y�$f�*���_d{�u^W��kǈ+�F�5/,�L�O�NhL�+�s�= ?q ѭ�� �b#ʳ�-aBw�����7h�B<��3)��!T��v|���M���B�П�ٗ	�>ڽF������`���~G�n��<`?�����r�����q,�����H�G�������w-����^ {���-x2��ez�3���)@U8=H8�%KZM�4K8��`6�X|�D� ܷ{��}�mqSj�9c�H@i��U.n�5�\� 5�1�
��ع3�<ee�3��K�������&�e(�AW���Z���L �+���O���@��w�ʔ{�R��+�X���S�ր)�:u
��t2��t���k�[�=O�&Q\n٬�6ʊ�85^)���^a^��V�!��Ә���什`�&~θ`:�<��M SO��|d�*;�U�L���0=~���O�� ���lﾹ�s��v�.�� �g-����{r!�@$�#6=]*v�a��r�e�jsX��,/O?!x�^\���Z��E�I&��x�Fp�������XB*��pboC�� _�\�a�!���K� Ӓ��#����7������3!z#�}�bsb"O �8?�ʞ�� �'M�Gm��݁�W�:���#w�DJ�����Q��s#E�J�2��M��L�۴
�$]^h���Lw?��-���=�+*<��K�Ud���y��XƔi�8���c;���r�o�:��J�O��m��4`I�
�ѹ����|��s""�: $�=f�Ӝ�fOﾘ��*Qu��k��ߜOrݫC�5GTW/ӆ��������^y��d�O�d�@�	�Oa:�y7�(��xޙ�O�A{��?:�3�幁k�l�����>)#�q�>���F9���I ��K^ם�^��B񮑲�[��^��2þ;����jgOCڑD����BHƪ:���4��2j�%K���J�Z�����Xp^�^f��u�������O�K�/Q�]�4ҽ��!�xӋXE�ր]�w��*�Z8K�\[�dN�#i��@�Z�'���J:1���3~�7����l0�E��2�1x�Ղ)��Xce���C����I���#IP�K�.6y�^�n��/i��L
���
�V�b�ҽ��������ZV7�.��w����/kO*�� #i$�r��x�M��b�ù��7ׯ���x�J/�VVQ�iDw6,}L$|k���#z��������,��ѣФ�s�r�:٠������_>����>5��� �	��T��}<j����X���U.��������7���x^�i�`FZS\��S���'�tc�Nins���e.������Dp�A(wy�is��l�p$��3=��8�� \U��������ޡn�9��
?<8�H�96��hW��$�"&�Lj丈;}Q�My�p�C�ZX�}���l���l)�tQ�pq���] 3�ݿ߲�4N�)ժ˘�P���>d{̻�����b�Ր���?Gy�[�]/0��tQ�H�r	�⯦QvRh�:I����F^ljF�-8�M�\L��j$e�ر���)������GW��az�H�ݓ�[y���T��O�!q�P�itE���)�D&�@���	n�����mu5&ɴ �tB��o�AA��B��T�0 ����O
��q�@�^�@�j�A�l�@3�?o�գ>i뾂vѣ�8��l�r��&�w��Μ5��x�m��z��n�>a�Em�lȹ�5�	CJ��+�O۪c�@F�Jԉf+��W
[}�������2�l .����H��~<R`>|��o��K���E\�֣)����U�V�]�ɺi��*���΍��Β�R�f��I���F�~�> Q�r97�a	J��q�8�Wgdʦ��-6@0~�0z�a��V��4J�"�1�A0�u���J��Y����^���u���&P#Fx�0���$��B��+�">����M��=�l�$�-$��2�L��V5���0��QbAIXҋ��vS0�U��`��ٯё
�
�F�!r���ʩc����h��LM1��{E�-�x�Su�Q�-g��T�r�|����j��<���]V���p ���'-�P�ˇ�f:����K�� �ӓ6}�9Vj3D���qU���s=[�3B�~��&	h�U��px\�d��+*[��QT1Y)��7of�8u�5�E��h��ک�ݥ�{��&"��'KEc�VT�N���F�v|��u�#�U���e錡_igCI�Dt�a�����iEn�LG��*��z�a]�D}��)r�S�ӯ��-JcPwF�,��{�Dr��A�[a���7 �
k����_+�O�A����v)qu�<pH7�Y{��ܩ�W�%�$�׶�_�(�ι�f�S$�N�[�[��u�)����Sʉ2�)p��hx�R�_'�^k���đ,�&�����N���kb���2�:�����3���J�}{u�ج5]#c�ѝ+D��#�5�d�$8���R���T2�cF�S�6�D!8,��A�w<�3X��	B�jE[+
]Z�WR[΍,}?*)��x֔����E�'
%)���S�z*��!G���=�@T��ٻK��=3J�+�9�"�,���*����
?Q�l�X�X����^?��aҚh9�#w��"���Z9�S[����:�%��Ys���5�Y���^P`e�Q����v��[Τ "�vV�C8<�!��7���g��
\��S)
.RF"�w�%�q���ڧ�8@�_k����<o���V>�X�ե�H$�0����P͘gfH�̍j#��a^%�2�K�Q�������Y0P��������ѡ[h�4&�I�i�u#Vf�
)FI���|p����C��m�w��@E4t���oD��,����p&�3��mn��muu'ٞ��'��iI���+g�ΕN6��R���`م WF�F��6|���d�۝�)��`��TYcDx*��]�����'R����]��nϹ��ZwG�!R�HY�h��(-���9|�4����j�]7r9�4�>��&�Ќ��4~.�Qg䖅�fX�ʞ 8�ަȆZۄ�w�?�9�-$�����s�!��)��9�o������tl��/�,�wv�Zpiv/,q⽖օ�6R�k :k6�D+�A�)�]��baL��]�-����L04��wvw��;M���q�0:@�dgahf��@�Vb�	�Ҟpɝ�SBв��W%�^ =Ԓ�8lr�Yq��k�%�.#������DN|�.�"�# ���2R�����#?ee_`��.U�L�1��Ė����Uwr�W��fI �	���[��/s��h�%�8?�]"Gؠ����l��������;�i��^ޣ>#(�9�(9n
��t����V�D}���mSy��[b(ƌlHB/ �N�b)zpxe�ơ�KS���#��L����"/�:�T�潧U��/y�(�^���57~9-����@Z��l$��e̔�F���~e���jS�8[bt�6۸.��M]��O@BK�����2(�}�<�I���djˡ�8Ҋ{юJ^��iѴb�k�4QTԧ)�Ms*�P�g%'��=9�=L��@.���-�Z������T}��8���]P��]U��N{GS�����l4Ka��Z2'fL3 {��e��_B���s���Ξ��[��͚58��*�[��P���
�F��N��� ���4ȹi_2��[\���I~�`�$-n�<���D�S��a�wk|
	|��s,:Za�1-���e�G+�`�an�;V���;gi��X��A��-���`&ث2Q}��ߢ��| +S�W�:��p!�#6���i��!ʘ/[I���*[H���ӑs@��ae1�\0�^�ਰ(�
Q��B�s*p)������L��&M���#Ooxt!�7�ˮ�{�;�}�4$=3���^M�o�چ�9��H�o��mY���`~ܤ�H!X
�F�D�˚;��<��$S �ܚv�d�t��t��_՜C� �ਝn;�����ale���k�GR��={��wc<83RP�����rg���QV�!�ۻV!��/2��X_)\��LW��R	&n!m�'N���Pv+�d�"P-���mi��������;7���9|�Z�]DH���S	È���<�{� ��,[�)%&1~N������X}�~"g�M��9���5JNx���(���`��D�U[J�W�������hֻ���d�GO��0�?�-��C|(0/c�X���U���*��>���Q��Cj(,V!���`��1�z84eW��e>)|���Bp6���&�3��b\%7�% ��
t��7�xi��۸5Y�p�!nF��ȷn`PiF��-����,N9��<�Z�C?�1|�v�J������2�#4e��h�5�:�&��9��T�1ꩶ=
c�*��Q��54�es�:�ΥSw�wQVl�v�� &M�h��Ӂ)X6{����J�!�.��>.L��ɣ���J^��������r�	z�y{���4ц��U<�����ĮV1�pTl��ev{}H������������0�\���
l�R�s� �[h��4a6Uƞ79�Q#+��*�W8���ۛ�z`L��o�5��L��~Zg��:��@��9���J:��s�/L��-*�|�3w\Ph�BP1s}@P��mY�զ�T�A�89z���?�\�n��� I�����&`��YV�Ey	�<:SzlI>�q��౪1^
������8w�;@�G�ԙ�u$�J1CT:�	�<����x�����(��\�����3#��Õ�՚��T�������r�l��KK�:�l
u����.��=	��ϼǄۓ`�K��Q���2=>Cpvԓ� :y��=�w"�ز����9%hᔕ��Y�tOI��
FN���ut<u;��F(BD���~بk5�qm]�2r�2����Q��+C�i�>�sCS�͇���[��Q�N-�1$��m��Ug��T��1�9GZ�j�gU+IR���ޝ���INF�%�χ2�b&�
]�X,���S� �7c<Ţ�9��U��?�~T��2�.�M6fe&������Y�v�)�K�.�zaM6Y��L��u3��|��N[�S�;1��4�(��#��E��	ק�ҵ��"휋?Y	Z���O :&ΐ��Ň_S-��h�: ����a���%3/H7W*��k�j��fjb�/%#�q�?ޅ3��M��.7;L��Y��hƈ)Q�|��*���}tBT&ꢔ��ML;����M��E#�lOH)��W4A" 8�2l��i��M�._�v������Hd��F�6B�h��9���l�bu�a(�p�b=&�i���d��y�9�ýB�I~Z:��9Eo�*�LT�_U�b�d!�Ü�V�@��=_�2����L����G ��5� `�(e�蘩�Ib%�	:)y'��a��b�pQq��DN�HS��ܕ��^аYˋ |���*�"�@۽��5pe�Xg�PI'x��`���u���D<�(�*)��D�����4����{G�U���t�m~J�J[y<�i�:i��n1��u o3fY���B��'o����C/f�-���yp���[� w�K��5�v���Bͩ��7+7���Q2��uH��i$�~��� �B}����M��,��E��M>��E(Z����W�k��9�o��Y)j^�v�BM���� -���a�-ql�k!Q�EL��w4C���=���5b�O�C䦛�5�qGԥ8w��^� _�� �j'�wʀ���ъz�Y��|��vl@���6>]�r˶��-3f悥�&kv�;�M#�A��U�}�h��n�0*S�75��j���''���H�a�C��U����~����7�����9X/��.^P�ܙ��(���u�P�Df �r�<	:D���n�n�
uGᏏ�
R�pd�4%R� �k�|�}Bcr6r���X�^L� �(�-mwܥ� ��޼'�m��:�tn8q�B8u���]�f.i1�$a���������#����;>��� �̞[c*f(�p"F�$?:��x����zv�!�V����b���UӨ���!�8�.^�Қ?���g�xl��?��?����Y�Cw�T���H���x�J9ώ�ͻ����q=Js̯Q���	U�G�ˬ0��V8Yҕ�E6{�9&Y��/���֌Pj�J�|S<e23jZ�J߀���ix��ik1X��#b����xB+@���*�Lv�����]'�5�<�C�F!`­�D]�_̔.7')*̡;���R�񨼆Щ A���^�7�Y�b����Ӱt��k�K���
�t¥ߥ���{Ni`��@��~��x�(?���-�@5�;���]��)�\��/�$�@7�v�~v�I>�.O~nK'��*����Y0�W�b2Ć���r<�8X�m���3n1�'�t&��Kg���B�C���,(���vf_GħZ(����_����AS����A��:�N�_<���j�j"�M=٪%Qq�텚M@FI�S2猷��9%��[�(16sW�vW�ڈl��hM�Wh��T�D�sR>:p*�f���+*D���I�4}�h�{�HBe�g�>���a���n�m�����Q:K�3tw���eT�g�W���}tm|D�H�LAsz��&�c)�&{�ZP���]����	Z_\��%8��������x���[�P����(\ݪg?�T�
i)�"C��61֑V��Wj�Xo�zO(����=�����%>��%%�7?٢��gV�Eڄ:>��tnB�.���rQHKlzh�k�"����-Ó�Vb�)�����@��$��ߖv�}~ʋ�	%Ғ�u�n�i8�7�`G~��-_4l�*���{�[n)��n�fiΨ?`l|�x�@K,�p�,� ��ڎ9�=yl����Ghr8��.����i��V����z!�`��b�TT���n�+{'��%]�mPx�L�����@����J~Y���5XNJ�__��DC�'ky>��W���
���m���S�:9����LI�����FE�FV������Va��"xܘ�����nz�W�>�����̹e�F�q%Y���s4��F5�Ӷ}����܌;B�f��O�D�7:Q)�e�$}Z�G�Ո���ǒ�]Q����0%)㔒A;b+��P::3�)'pl����l&��?����EG������Q�A�cs��(�(���9(P=������8�R�7�nXjYi��T��۹���0����d�G-��4����� ��WGhM��՛���aN��?�H���q N�m��|���d���g(.Pе���yGa�I���0�$��iy��J��(nI��2�1ܷ����l��,KZ�RZHYa)!9��3�dd� 8$�\0�����6�.} [07Ɨ�S\/����]פ�>?� &�`OP.�4�Z]��BD�����bl։��κ��tb�����{�g�/�"(�4r�8A:�P� E��[�9�*����Ѐ]ʨ:7���M���[���/��g�Fm���5B����8��	\ں��^D����=-T%�caR���������U�	�H��SH�ŵ�H ��k>����qVM�}c]��_��䶑�tF�&����"�LL��8t�|wyBq2�C�ހ=Y׋�Vd�hz���J/ >�>������ʤ��z���J3���|$EXJȁCEW�B����w�����,�P�]y��e;/
��ע ��u�����K�Co}��z"��3U�L�?s��f�'yM�䖺�'k�wS�2��ԃ*�C��4�^y�>���^��G>�����NjNIB^%<�r�f}�k�-Ð{��8qi���x�ggR�܀Q��Υ����r꿾�_�	�<��9�������^4A���X�5���ܕ�԰'b`q��b�* ��v��2�qJ��Y�BϘ�:³�%�ǳ��A��#*7�X�w�2nȝ�+F&�夔�Mb�X��ѣ���d{�hٰ?�[{�����7�:G!�uv��	H���p����8�/h��3֐L���.sH%t�=a;����\^�B���.�nyz;�.T[b�����m�t���ٜ���j��H��[�&�^�Εi�so����DOj�������lI�au����U���b�u�׊����-J�L��8�lѵ% K��nᄅ��1�,ZH���Vn�SU4\��Piv�MG
����g��� �1�!����A�7��t��g�j�`�S)���/���#`ѳ��7T����C�u7����<�oV�
#�L�ol6r�TXI�z�]����rr��������HNY�䜒
8Q��f�B���F�ˆ��5��Q�wOE
��w��yk
Q.L�>+��D8�~	��xNcF�2?�ֆ��Y/rS���"J�N�.^#�*��j�l��oV`:�B����fC�zl�69�p�(ك)�U^ �$թz`}�͆��cu�Kl#V�Qdyް� ���%.5\�>�|�R��L<]�+<HqE�s���e�d3��њw�Ok�)�X��xt���_�����?5�\��9-Q�z(%���g���D�����қ����(Vl�{�>b8J�}���;�����d�e^�g֌3����)�Sp�T���@]�q\��K���(�f[���r��o��^�S�nhr�V$�9䶄��;� ��W���W�؞xA�Y��h�3ENg��$�_'�u��C�pXNEA8�'�f��E/��}��8��a"/R��G6�cw
�n5��n�F�i�m��:Eue��g���uA]FD�z���=M�ƛ��B]Z�Sŀ����oA2�����:�	pd�/C�'3+��Ҹ��nk�G]��.�a�кII#�v�^�[O�>��R'��Z"���U'!�[�D��,J�rS>��s	I���2���/뢿8N"��B��������2�8�Q�\�v��?;G��uC5Q����s>np���-�^��.�����74[��D�q������	Ư��k<��y�e�V����q�A\ R���h�hT�\��k��j��������n%i��zU���W�*hC�H��+�s���N	�ܚw�n؍�|���|GF!ӁS����)�aN총H��2�<��!���߾���I��,8@ K��r�i���M����ջ��X���*�h��*g~ "�}�d��e����'5�Қk�z�2l�� zFL�e��&$��Vf)�>E��w���w�#+�����h��R�w��f^qw�9��ͤWN�vH?+6���t�W������p���Ա&*ޓ�ٿI�'N�R��+����X��-������w\��7k�{�W��	�A�L�g짦;�K�t�sg�Q���ϧ�{�M�9�P��a8*���N��rc��]쒚7�I�������Oؐ�bd>���練�� 6@��[�.��U�F�I�3���e`s̓A��=�@Ց����:�i�a8�u������2��=�'�2^����"�+$��r&�N�r`Ǧ�qR0�pv����	e]nJ-*;<*������b�P���45zB)3/G���ui�Ifq���X`�(E�6@�j&q���VQ�M��,�P�p����zw������&�|�8��8w���㶻� Ub9�%Yqi�$�������S28��+��h*> �TƮ�Λ�e�f:`��x����Km�j-G����� �"F�A�Ќ�T��y
>l�h∸vE����#Ss��I��D�&ɡ�����dӕ�}��G� ��<��mV�iİ�^~�v0��k�W(���!"�.M=CH.����[����������KW�g�{#�h�w{��"F� �
bn�Ѻ�r�8����hj�;�%��2?K�h-R�H#o���C) R�B$�{�E�r�����7��af�����R�e�8��/0G?��Ӫ����3/U]5lt��.��@�bE-=D��)���7��u�1mՖ�fw���4��ם�����X�9�3��K�2j!���A�$D{\3:�j-�u~M�J"SV��ؖ[gx����\��'n~���2��:9��/n������C���S�D�R5�����h�q�o�6���/u���K;���ih#��ȓ��WW��]܄�ܟ7j�6�B�Y�҈���%��B=�}s�(t��ҭWޭ�M.V�?w@�����m4TTҭ�I�s����%,�y]��<F��h�ڇ�|��� �ѕ�ʥ2��T]9!�����R8����K���fZ��D4�О6�UA���(��ʥt�,'��mu�ޘz���{\JP[��@<o�Cۮ��0{h������N�k�Bo�?�r�˯!��r�d�ti���j�2�{�RE`h�����2�[1��k�S����f�M�tT:[o�^V�\��x^��A�����P�t+O:c}k9���3�&�Ur���&ٷ�#s`���.�	>e�7���g�S��h ���w����gK��^��2`r+jW�Bɠ{ڊ8aoL9��g�@���@��d�+��^̆\iEN��.c�@'D�,3��935��r"tIN�����BzS���"S{ͷs6�K���P��g�?ݛ���F�8y7�Z�q�j_�+Z��tZ/�CP�j�}�f��L��_��:]���;�b���T�9��v�%�w,?wC@�������+��_k���:J˘]���*t�T�Z���Z��t�D���&�y�����?�t,�j�R��R���j����Ç[��A��O+�Ψ+�Yt����2�hm�V�C�s�X���=�ϵ�RD^�3MVF3���d�MK����2�#��	��upj����1d���|�� �@���	�0 `�����E�m�vHӵ��{����w����}�J��^PZT�>����mл�a���y4�>k����g�4!���|�D(W��֐V�y,}c��yq�k�d��3x�zz�S�e��~` �2X�m3њH�Hcܕ�bu!ҍ,8²/����g��dx4bCx���q2F�9�"��B�en0B�����	!���MZ���etF�̣��D���LH�Bǹ�I�MJ���0<�IJ��h��+�� :��24`�_�/@��`��)�<[����ƻ�	����Qs�?di��v�dI�����v�0>��*�(�,��hs�#~B�k�~%�3�b��
�"�e�#	 �[�o�~}=���mfl��|��{�smLBΠ��k�lOl�d�)^�l�]s�U���C ��Pvܪg��L��y�INt�������Z��,���V5i�U{�y��F��s�|S� ��2�xq���� 4�"��d�I�0�������S��^h��A����������f�L�=�1-��� .G���5s�Lާ�%��cI\� y�މC��V��0�>}�w���mb�������thm��`�)��s�ϩ��h�눢x��Q�+Z�ۜ�nX�ȣS�6h/qٯ��� ��B��Z������{�(��z��*`д��.Ό���v*:rRوs���ɷ�(��/��)՛)��>'��3�2��b�F3᳎��-�_��H�w�-�	mfY�� j����b9��_��+�io
()e��*r��4^�� <| ���i�Y����6��M��ʲ6L�I ,��y����[��![ϻ�pd%��g���_N8��.�0�ӡx/	�hֈN�=2�\�&���\J����-be�Z��x���BuD���h���Whr�n�;8��L�X�>���"��̾�N#Տ�1�\��>%�Cx_S��db�0�䪁"C��#�6)HOM��20p����? Ezeԭ���cw�'P@�Ͼ����ED��~�H�4Ҙ��h⍋�����7�#Z4PN��|�����L�e۩��k�J�'9�s��
�U��3f�dKL���%����[�؜��,�h^EIW$C�%�7c���OY93者rA��ʢ	���t�����F�����ء�5@#�d�l���d%�_n�x]�GGP�K�DN{��������2�o?T�����ԤcT	-O��#i�@���|7봷�)S3�g�M�C�F:���Cubj����	q��rR�&m�J�H?��}�{��W0���gr���[4�����L"s��Mi������m�%��)G�zy��;��� /�uВ�^�Bn���U\H�廷�pl�|��Uc> 3�Hs��K�Wm��᢯~�0*����{;(>���k�Hΐ��l9bF��|�*���˚�.�k5B�Z��TB����T&L*�W��t�\n�4�[�N���z@ff�������#���M_�$T�얚�4��˩6)掭���,�YƠ�A�dZD>��,ŒR���Ђ3D��F�x�2A�-�B<�P3}�S,"4q_Lo�(��r�T�c�vЯU[��Um�q�,T	s�]�w�/��,�S���YH[�kd������^��K���k�l;��)q/jW�O��i�C�'I��%H��F�Q�0k},س�.��[;(���V�����)�V���Y�j+��Z��9ώ*CX�>�h4�I��}	���^)i�@��),��n�ao/�<X(�PQ�u���>��R?�k�;3��4��S^Wh5��z��}0��h����6}��Ĩ6��&�K�%���-kQ������9$Py!m��Б.�Ǔ��+�0�a��%v��y����Fla��p헆���p,?_���S��&�yM�������!B���0�����M8�W��p��uW"������Ѷo`���g-j��0;z$d&��Wzا3�3Tպ�~��@�ֳ�RK��
���4LE�Uߔ����z�TG��˲'�?o�z���{�Δ�� ,DhiMʕܽ��m&-R �i����&�ܓC���DfN�����7F�������
1HZ �7��7��
��3��h�u��yA|�B`X_����ƺ�$߲�z��"sҟ(O���|e���._g^ȾzKv�0��>2Tƒ��o;�M ���
~���`N��w n L�F^MQ��!ڊ�F���۾�ᐣa T_�����/=?���)���*̆���c��<�e�N��FӚ��BS��|n����ë4�)'inT�IXi�m��=/�����ϓ`��@�	u΁����Ĵ���,.�_�T]-@�����-f���<����8�+iuV�J"�����T����(��ޚ��<�g��`=:�)�"���X�:���F�s�艂^!5~MB���Ҥ���V��t'���cr��+��5��5��#�wL��(��\�%G16`�եp30�%0���Y#Y�#��ʅ�}-�]F7H�_�g�c�lA<�̇�I���>*Z�A��hisv�R��m�[$1G�~o>�^�Аע3���@�!�4�%�����>;�<���貘?��ؤ�=%M�=s��nmC�]�/� j��Xe�uCg��0��P��`�ɺ�۷T��iF��3��.v���j�_���` ���U����}̋�źu%�H��Q�4�j�/� 	ZNP#�X���I�V 	`r�aI���Nehz�O�Ś�������XTu�9���c%��R�n�B�c�H����a�>Ǧ̈́�����p̾m��}�E/0#!��A̤�S)x>&<H6m�2��I[MT��;v��MY���bѢ��OsQr���s���(�`�|�ͽ�Y�a<�
�����Ӥ%������ȼk��iqԎ��7f�x�P���,_�:�u7�NR�􍁘��{��~�z`�s�5柘N�3��?�ϫ�ڷ�;l&���8s�)�@� �۠߿׽�dt� �h�S)�� ̊߂�w��@�_�#̜L_v�J,'�-n�j�os?M��k]�����#��	Spa"�e�{F�A<������~/��m��3Oʉ���s�	���"��h�:N�>.!���J �9v�]�� $����*���(s̨x18���U�.�r.#-s}�0�1J��͒��+��W0�WA��ԯ�Þ3ĎiqIL��g��?kTX�oܣ�k@�A�dJ�95{L��^e<���*��(D��&�$�p���]�1���o	+wl��d-�Q�K�Q�Z���u���X��NPN<l������p;��.=�E��#�+�o�.�� ��G=b�E���_椣�0Μ�I/:�L�N`b��T�)N�e�ۭ�D����D��vJ3%�ƓS�q*c��XW@ʕy�ݍ�<�X���k����Ox���������Ld�G��w�� ɾ	�cu1��4Dk԰��7}'Tg��c�Э0yF}N R/A�b����э��nu�4�a�eB&wK{�$G�jX�1������T:����UZ&3d�Y2��3׍��r�2l�ұ�k:�qT��@����1n�8�T��%?������6/�v=]=�wA�@�������w�T>��{Kk���O{�C�{֘JG�۟��C�fQ��Tq��O�j��}�֙H s�ج�s�5W3"t��O��xJ���s
�ׁv/��7,�K}�n�
O��kǨĲ�ZY,c�4�F����%�ǽ�\=ax�8{l��P���G{_��t:��]	��7�L׳���U��4��_���??9*YBű�l��|6���*9�Q��7$�r��k�p��qlb���]��}s�V��	Bߘ�E��B �%H���Z�ʽ/RB( �s��p�R�VR�S�+εau�RM��"�L~,���B�M{�;+����Z�7�8���D>P������@i�oV�_��OK󣑒��Z�Ǭu��Є���{�/>#�;��<�K�	��ͦF��1�����,f~���#Z��[Fvd�Rx9��g>�s>���)_Pw�z�����tj��Ҳb��p\�I ������s*;fyə�Zx$OGj�*>�`
�~��됯\�np��2}��K��C��v��6����,��Ox�Zv����������U��e*��Zi�َr��&�������-�$����
���\�ѺNך�Ԩ)(OA��3�^�Iɺ"��SQ�/�S�������H�9��۸y$"bHgz�G��� }3�1"v�=�%�K�wR�n�����!u�e�3gF���Zp�̊$�{���jCΦ\��L����֑i��U	L��l�W�U:Z|�d^��t@@�~����HLp�n�~a^ȴ7m��h+�65Я�l]ƽl����?N)���6y�S�w2瘂Mhw
��3_x�WLX�����sY�3�S�Ҫ3cP�t�;;N4�0�%�_�EbC����	�2ג���C*�P^���ih��q��c0��g�T%ǰ|LgZ��k�H,v�AU�h[lIz�<�3��d�[u�GrJ"�(�rIOէ?����rl�m��!yI\�"
����yсJ߫����%�Iq�ɴ�Q�aǫ8)�B�=�5C��U=���� ��f����x��1��ٔ�v|��]H+D�����V��Nk���eu��p��n3*�q�L��p�n���̈́�􊻍6W	�$���H�w��,,q�9���~��eg_�P���J�B�]jR��x�>W �Z���Lz������}g ���3��a�¦�i�@v�Z[�;+�Y�ֆ�3�r�ց��u��ti��G���+6����i쉯o'��d����'�f.��6�J$D��40k���ូX$�0�e)����t4�;��s݀�����2C��L_�}��s����q�=�����M�V,t�r�v������l�X�E9K��EF�u:�6&"���9�%Ƚd?�D< w2���(�z>�؍M�S_U�C�aT������<e�O"���B��`z@!�5���q­�3_�m1)�ku�$�j��(�/y�S��9��|T��cZ�������_DG�$C|�酉0 h#�JZ%T騦2��-�"m7��U��<�H��j����>�Slq��7����A;���vf�)�<�7��-<S�T���˺N��`�<?���V/��f#��u��Ob~m�->�Rt� �n��$�ƘW્o�x��4��Vȕ��j�ۨ����''�;uJ���-1�f_��yV����Ov�$X�� ��;���՚#����x�3���>��7D>kƊ?,=�|9�ٽ��� ��H�>�u[!FLje�-�R8�:��[pv��M��5�e�JD45�#�#y@�����k1�+�V���͑*��?Bv.:)nI���&��?	j���̶���#P�V{�x��©�4��tWmOx,�����OX"kK��nX}ݑ	�-�g�#JU�Sv�ﲄ��ʑQ)��U�E��f�߽��}�K=U�`�[ ;���wk(���*��^y~5% `aB>��8<QUy��'��T�l�i2N��T~ � �LM�DϮ1�Y�d>��C��Rh � �B(h���A#j�b���p�B�`	����Ͽ�L1�g���$�O��Ub����{�d�M�������E�ś>�]���6����,�0�~5������a�AHH�q��� �s��r�k�A\<B�B����Ԉi3������T$���d��/-a�֟����"NT<Hk�mJk3��2_�'}��`m��-��
�4�p���������"Q��P#	�!G��g�!5Hd�4�n ���[�%��u"E��z��!�-������c�-��� ��յ"�a|�a�	�0���쵴�;r������ �yn�5.�����9�Hٝ ��m�39�*�p�2��~_Z�DLQ< K�'�W�,���Ζ)��i�`�t�$�o��6��4Q�ԉ �i}�fvTg3+ҏ��� �dx ��^�w��p�!��'�Hwֱ��t�P��J��$i�ʓ|&��7Nzy�n^R5���8q�g���Vo�e���&�,s[�G6�T���?S��3*�7%&�s���� �4�[Jv��X��p��<¨�W������F�)�Fx�*4�%�
�]�����z�� 뎕lӣ�oB�׆��Ni�4]��qs�)ԭ�J��2��)��K�xܤ�~��틌>�0_������}�`��O�.��K6#��(	����*bu�ƨyq�>���O׶̣��8�����n��W�Te!7o:V+=6r�?�(B�ݯu Toh)���;�v�-j8}����Z#�����τۤ�i��X�y�;��̖^����'�jݲ��Ȏq�r�O0V��x�����M#�3◢��n�]N�0��p',���$�=�����G4�Oq9��X���VR�z��[#�� N��ۘnC�
��8EӶȭgMM�f��n[�����r9	� �/H0V��R,嗅���'ca�h��E�f�X#������tgn�r��
�տ��Go$>�������5�v��Q枩	�O�[&��St�qŨW��R��[���P��g>'|�-.�_�=M3�Ǔ�(������g���U�pdo�+,y&P��?�c;��M?�&bձ��%?"����[��7,? �i@�^�6ll����%o��	�@Q��Q��L�)��6{�$���>:��P)=����F��jz��)�4'�*�`f^��'B�<�`�G�xп��*�?��K���IS�zy������'���Zh�����c���89���j�L=��Q�F�31���V�:*��R��4��q�vnUl��L2c�1�0&w�H��B��2g��F<-��"b�Gb���J�&L��\��VIhѼ�ª��ۇ�(m&����3��+�V@�tY�S<�����6H]mu�5s�9�k-P��I�V� y�}�{��!χ�
�K��H�V�A��~��,��ݮ���	Wa�O�ğ���e֨��Re��5�.����������%wm�J`�!	i����f1�m
	a)$��Z6zw��Z l�IwF�"���ѻ3�sn!�'u�A;��̈́���V��^=0�}%���6�k�1տ�s;D
�_�8:M����gY�';�<o�7ڌ�"�[���k���/�4=�1i��C�}��8;�8|®���:K^Y�8�ǹ�d���+�[r��`w�z���φ	R�Pp|�L��amljaݺH���@f�@���]E�P;ت}���}"1��ٸ~�dL@¹����_x��0ö�Q_E�a���<����S%V{c2����]5��8���g[H���o2����0�}xb�X8@.m�d? ��aOӗ�C)1t�T�S�|m¾�F���UC���_�P��}T���=��Ecɝ���Ρ)�% �Ķ?�_�m:j�=_=���F���i6>�d*G���Nӟ��t�N$Z�)TT� (A�$#Y<�����+ ��~yM�*��b�#c:7(&g��*��@o\�B�):~o�h7T2�R:E>��
���7�H�l5��Vi�T�J��$Lg�A����6�~,�Lk�̽�ٿ��7���ɛ��Yp �_?�e��h2�?hhҴ�Z0Ki� B�=GWRۡ��A��Tt�j�zk��=O`�ϳ@?�E�N�}^IzN�cnȧ�9��u�fCoRQq�V8�m�N����G9>���Ȑ�M�v70b'zi`䬞QG�fHiE.������W�03����������[����}4���e1P�6�'��xKE�6_X��ME[ʿ�Q��0��ə���-����eF����{N��Oe�it�K�:�C�����f��\`%{����E�">܊�y��	^�l1}qC��u����� ���&�R��M�ؖ�p�g.��K�66��1��B �;S�g��k���nI�Ѝ���V��)z5vY��,���1F	OCX��B�c���!�~����J�PjA�XX�?�������]Y�_�8�i�)�>�o}P�ck�w�1V)ȳ�C�k◾����U���b*i��3Z@ý7��ݱ��`�S�\�B	!B`�������jT%�>Q��'��!*�k;� �P�_��s�b��d\����0޺T�T"���b|�������
�
��	����]m�ݖ4_P#V�
:�L|�ehP_nژ9}Nczw����U�l�d�&���-��ÐEM�Uɒ�i����u��a�;�t�pS҅(�ظ�ȖH�3̚�Gw'���!G�c��٪�'�I>ul��M
G��%�o�<NUީ��}�h���eQ͐F��iY�ptv�FFP9����^�&�(� ">�.HZ�9\J;�)�2ԉ1��y�'�\O���)��tC�2x��;�5��;�LZ�sĜCj����{�KI=8
 ��i_��?u	^�T��1B�g�^D��}KTl8�f�P/PU8L/��Y�
b׼���Y�zP�\qI�h�!�4�+��Ȫ'T+�@p6�`f[�b�֕%��0��6M�ص=@����GMg�)�*��ȥ�E�l�_��1�/�~c�~L	��V���EQ�K�h�lӇ4e��E�O{G5�M�E)ʞ[YV�^W�@�
q��@j�����Q�^tO޹��`3�&��H�B�<�fJ�YS��I�7�Mj~��D��'M���(�m�d{K��v��� ���,�>��sQmf��U���F������:D�xY`d�H��$�+Y��C�{�����#�t{"D��ʾ�A2���-�<Uv�Ƴ�����>w��L�h#�+IKV��-�{�>�~�y�|��H�����iL۪�8��[y��9ڛ|�pH����}py�"�E*��?�k#o$H6��6�����f�I�?J�B����?�'���c���έ�{��=��Ҁ+��ll��h_��X�
���ٌ�v+�&�PɯZ�������in�a���^UB��X�ѵ$��Nk\Pk8�T���U�,
$a%a1��$Ws�m=��ǘ`�ܹ��dcd��������?�"mm�VrIFÏ��sԃ�ĝ��r89��z0�E�]��Ef�o���os��'3|�F$�����4��d��&2.���f<-�՚��C��g��('�7>ic��}�0&��H��0&G����3E���DԞ�3����S��@ǣ��ٻ�d����$�̹N0���T�e-�O	����F߮��]`Ό$�~�R]�,-����9�y6m���7����y�a}��$�(���>���("r�t��ø�e�<z��/g�Ć� ��h��?�o��Yf��`�|0r�
�w3��Rw8Km�ni�ڴ��2ܫ�)�F� �K3!�,���m'�� �mVR
0��g�]~���U�1B*�s���EQ	E3/侍�gM���|�U+ɶ��;g+u&ӈ@���	#~��Gd�*��.zM/mF�т7h����C�#��?8��蚡٫��C�pZ>�/亵��4��n�������c��T�q�	~8s�Ć�զ�<��k�m~#\��4��M��֨�R�Dz�*���CT�gh���Г+��$�SEC���d���y�(���g�mgTY������d��ٺ�䀸�e�4�;n�!�k��Y�T��|X=���}���P��&��k�����xu���rڎ;�[u���������.N��]iذ�H��ThB�
#K�k����ƈ��38v����s4��[`5j��Z�#c��D�uQ�"��U���Z�ʘde��N,��[��bj~D�G 6�ב�WL���@�9�C�+���U|�d�B/���H@8�Y��w��a]�[9���7ʧ�
�ٍ^�8
0��׽pO��E��	\~IaՀ��ȟn"�lk(�Bʟ���]�z+e@[����\�ߤ�9N���8��Y�q{���Nt��_�B�j-J�ni�M��4]��}���e��m*6ȍ�|8���璳�8q�X!�����Xg�Ҥo�5ږ��A�P�`���3�E=�D�Ȗ�E�0��|�%���?�B~R�埜��M� �W�n$*8/����	bj�n�>�zs��Y���QHC@��(?�L�������>I��n�Cl��v@$��2n%#�۰�����0���rU݆�>����A���^_h�
�e�P��	��2}�W!Vo�g����2A�1�2bw���Mȓ�\lm�� �
Qv�2S�P�*&�����,y����?Fd]Q����Ss|u)�C	�?��{��ԃ��M�Q=�ν�V����^�|��Н�-dMxx�-s<�&��ƺKd׉�ᓨ��_���Ԡ8ﾨ�I#�fDP4��`�Wt��p����|,R���Ga�~3�j"/���A�3��E�m��G	`���ˊT!��h`�$����T�2�V����`sa�`1r�mis�إ�v��_J��}Ѻ�&}�{�M��7��olNz_��#�<�W�邸��ڠ��@~���C�M2^��%��rK��mB$� .��� i��C*����-���Ԃ�Lp-mt�t��N%XN�v=&�O�ө��s�g�0t�',�by]�u� �P��8�v������y�����A�h�=�%�ڽ"������6S]hKv~}6�
e��6��j�X�e�!�҉����Áϯ�,�T�b���nV1�Tl�<!�|�1�(R�-���G׳�\n�H^��:gc���x�/;�h9�?#�P�bu�3Jx��$��[=J�5êU�U蝍�Ǒ��O�z���1%:�r����-G�xU@��-�w|���_W���]�75��f���ʼ�cj,�
��V��;fgﱗ%��9O�fH]>Qg�0Y�r���-"�笕�s��cZ���Q:�{�yp�< ��9�e���T��~]��SXrv^�Ӱ�錉�f��e���	� f*��r���l������A��5X��#>h�L�zv%�.�U�
��˘J�\\�b�����.V��[��ع����bP�P�'�6$�@�d��L��`pT��s�Y1v������=w3��A7&�j�8�&�/1=��DJIAƸ0���K��3���9j]�����-��c2Н��g:�����=�W��c��fß�6%.{=>����H		dd|Xh�zN%#[{���`x�K��+�d�+D���v�Vħ���ݽτD��{�3SLfT?�j�w��@>o�c�u�o�N(7C���ݍ9�buh��z�ȓ�V�]�9Stw�+������\-������ک�@��(�M����ɤ��/�w�/ti_��;�rw��-b���E�֙��Š�ﵒ��ҪO	���{�hSa���F@�Xc;P�8z�<d�G�9t]۳Pr�������'����"�*p���q];��2�ǌ���i��G��p�NL�,�O��tqv�2����ːbw��Ƭ__G�r\yn����t�7}1������3Q�gz8�`n1c2��ZpB;�$���bl;E/4�F�/���iK@�8���냠c����$"�#�~3��2�7�(��rI��jnq�Ҿ=�.��������ә���LٰdO�sS��sy�d�v:p����n-55/�bFߥ�RC�A��Q��� ��F6�zC<e�/�^�P�h�����9w���<�h�] p��"�P�4�4<m�Z F�+�{*�a�5*�=��� � s��788.��X�|U��z�^~hOw
>i���K\-��u�,��#B w�9�Y(��w/cYK\fW5'b�$6�\�4���G�	 �)l'���3��u���� ���������>Oj���5�AY�<�Q��k ��b0H
;��1e�/stG�����0��.�/��3�:�
MP%��`|��3���<u�C�-� �N��W0�w���6���TZPp�N��S1�id�.�X�N F�%�Cz2.٧>1w���{�/K�.��)�5�C*||�y탑�}�!���jB
��Ӑu(?]�s��q�������i�~����t�j�`���,FhW��X�ӜD�!�l�Ϙ������eH�G_�1qSȄx>�P�.��AT94jB �7U�a{m��A�����ݔ|�ǅ�J/J?��x��ז�v��'e��	4*9���x�é9�*����q[��^�8x��T��q�G����8��� ���y���B�����h�9[>cJ���Baa��?!�]�Nc���;�W��6O@����o_���\�mʅ�=<D�_K1m��+�n�x��	;���#4p���� ����ʎ��Ʈ�[<o[������U�ݛg.~�%����Y�B"_՝�"�o�Z_�8���Hc��9�\� �^]r�.Fp���R�ܙi�V���td\A�e�o��������^���5�g��ф��z�� Q��\Y�k>�=Iw�d8��S ��礗���1��*�9����28��߰wodP^�k�"�m�Xq?9G�UW�S))��\By'�n��%:�8�"k�9�-��<|�0$
����Y�t�jA��RٝA�-�hӰ�w����+O�ue��</�史O1x�j)���O��uQ���h�N�p�Ɗ�%� �+�����j[w|og�KwR޳���~N��V����'��@������o�gИ3�X\��y�R�~[H��A?�<���녴�W8kQuHٰ�}�"LфvF؜�񛧆X}���[��6C �ބ�2���=��5����m�E,�mT�$�PV���r�e3���e��C�[{�3x3,�ۋ��6�M�*�8�7�]g�������r���K���0�O�AA�����>�>C��M�5(΂E�i�a�]�iA�+��T1 �"%��)�ȉ�&��q�:F��#�v��|aA;������_#��-�T;̺�P���MEq.R�nUH�J@�����<"'~HP���m����}q��$�DZ����e1���u�g���G``�&���>���p���Ǌ�0|7q��e�Ni��� ��ǃi�\-�Ƀ��(q2ǫ`�V��u�4(�7l�ft��5d2��
:'�bM�!�!�l��=$�0�U�!
�OW���߀t ��堂H{�g����яj�ۚ�����f�o��,���Y���t,�����D͕|[��3q��qݜtg@Z�����#;7���OD56�W��
z2_L4�1�/"Y|�Ieþdg���;Ҹ9풞)]^���4##	�QC]����7�EmP���%�bK<=wե��u\6ߪ�1�-��.`��0r����dH�&,T��C@<��qOf"ز_\7d2|$c�����/$	L�t,�c?(��ۊ��i�uR�i�Bv�
�-dȐ`%���\Ή=;�К0:�dk8�J�}��5��� �i
�D�D��_-��W�YD�k�z0�A=�-g��A�	{�T���pc%ט/�O�����'�_�D\&�yW׆��c�P��W����F��VFQ�s��e�&�N:W�z�w�����>;�Y;�v�"�㋙W���>B�:�4#q=Q�3�o�[7�[n
U]�A��F�Y��3��g]�¼$A)c_��� ��̥��F�?�d�84�r���k�b://Y2����}h�D��e��U�$ps��+�c��s�__���N{5�����t���d�݇��e^��v��D=R��:M���b�jz�q���P5^����Q0	�̘��_�<�.+����4�R�u�=�{"�#D��Dx��.zӇ��Xq�d�m*ܑ�ր'�j��
Z\:�}yJ�\u#Qe�� ��j���\Ĭ�u��y�h��D���ɘ�s/J�yr�T�PZI�F^��1�Ič�Q����\Y ��//@6R��]nZ1�wm�w��Z	�Ъ�{!4_�pK��n���3Z'e
��R ���-·�/BA���b���o�������$�?�2%��OC	Z�qn���7�J�ݫ��Ӆ	6"K��~
b2�E����.*�M�Q�P�x���L�Y͉ܜ�+%-��ґq ���toa��' -�+voX��g�����j(�kh�	��n�Xvh4`Y�o!�}��w$��t۰ �0%T!�\hF��{��BΝc�ԗ߇�2s}��G�n}O�����u��N�%�O�(�b\�w�a8���Ge�r*&T��
�	v?՞��סU��X�$���D�i�N����⌿r��G5��X�tk�v�#��>C_c��b�H�5�Zz{�Z�ZL��<3��l�2��|%Ҟ�k��ޘ��GCR�X4$ՙ1���OtT�-M�%�#g�	`,�A�N�.d�Awk&tt���p���"l� �f�D���RK�5�����kCo��aPH��@-�:M"������wF�u�G3믋zU$'��>�IcU�3�M��DN�UPK[��G�&^׶`�9v�έM��[9[��t�q��0�Y��;7{������U�Eh��ϥ onXB(���M�y	܆e�b#T&̔-���ڵ 3��.�n�� �\d��|R�����X1�d���^ꊤ/�_<d{un���bL#~�|�4��2u��i�ˈH���ߚ?ڨo��݂�_��<Q��bG� ma`-!�=.�!JlL+1��<tr���k�*x�[����c�(,�-�V{���i�m	�(X��!/pu�'��qJm�ր����w`Uy�O��@ͥ[,��f��K������ܧ�����=���a2 E��1�S�'�b0��M�0�(�EE�E������d�ȏ���T2j�aWi������]��l�F�G�����I)Pm�`k��>W>m܅ԗ����*u��4:�����Oy٣x_VZ�;j��{ݎ��p��]Ǜ���0�a�^,5�ض�5����=�<���}*�&r$�A���vK׻�����q�O���s �
��G���޹ *���_��#7C��La�%�T�����_ZR�O��t)�y�.piD�A=������`�Z���+���/X�����`�^�k�Tf�����g��[	�EO���â�<�I��Pw�ε��m[���;QU'l�T�M$m���W�� �`oDy�0y(+�<3���[,��ㆾG[:0	ȷE�mi�:�%�M`U�n�D�b�'̻OT�=��%>4
�X�ZߖI�f,����M
�Jf�)�E�m��I��5��D�kq�!Z"�DfzH+
�����
�-�9v��# �䠏{�l���p=�@�*9Wvz��5��$���
:����:=mpis�56����2��t�g�G�d�F�e�3��U���s!�j]z�;��[�Mw=fy�_,:0Rg%�vk�f�3�̋�}������es!g8�½
<�6��j��ÕZ�`�H��v�Ch�iu�/�D^�mHs(V�zشM�����q'y�*{������T�s�@�T�wB��/uJ*2���m��H��j�����?���A`J)�[�U&(�)��l�L�3�E�Ka�9��̑i|�<��r�V��ku�^!��	�<H�>/���Z7�Ç6mQ�}�x-�]K�R9ߜ(�C���5�q{�ZP�#�Q6N��<16h�F�g���� �O+T�Д�!�DCm�'"���N�z�(�BM�x�.Y�gX+zW2LF�A)�Q��s?��fx�˿�4�王ڛM��Ԅ|�T��Lm{*h�M�;:XM!K�2)ѱ��At���N���n����T��9��.h7J�I,~/6e�r���{ֳ��P�!k�!\-l42�,�c������� ��|hW���A�6�J�Aɒ��|�N[��<ﻨ�
�J���L6�{ـ��ӽ���/�]���	Wr��s�_yz����OOp�V��O��Q�C�7=��)W��_>��}yՑl�4���h�7�����E��G�dV_�y����@8=��`��I����n(z��iq$�t�4!�_%����7����S����t�v
���r2� �V��D�K���;aqjry?�=z�������oĎ�R�\���K�����U��j%,6�門�n�&��n�9�"���.q�ʵ�i�Ĉ&UW]���[Dћ]O?۫u������̐&�	�e೙���7���b�� �n�u��G[P�;�(y�vr ��c���Ct.��ޞ��)�T�v����==#7F�����'�n╇P���5ùöojC�M׋���u9����N���2���s�$Ԛ����5������紡2�H�wp��#��-,�����.��t'?(�:�T���-�λO���Z.\&Ic���:����ޤ�_mS�4A��"C�ݏ���5U�r�HAՈW}�"�P�w��TH�)�;nUJ���-�� ��}j׌��H�����X����6��IwDى�.Rubl�`f��0���E��%�{/Q"^�sN�rC$��B�{+)�Or#������r�E������T� ���-h��>d����-��8˶��2��Ͻ�D�cރ?ld��c�,�À%����^��2������5�hܣG�ܳr��.��̐��y�H��})�!KP�������x7�1�cY��|����\�ze��,���.��&
GP��T�~"1Eך)�G'�����W������P�

�y����Fj�1e�iX�m+�T������<�L.;�y��;���=�������aX;�b�X�L��RF�$U5-������Fb��Ao���{�.*k���@\�ޒ;��hmu�)<*V7pҚ�b
��ȓ��+�/?������d���00���R�� ��� H6Y���uK�C����S���HŤ�L���N����Af��q�����u�mt�;�A�-/-�N+6�#��j��HG�T���L1b�G`C�%�Dcz��s���\:�pY{�/a�N�5z�<Hy\m.�ykA��z�3�Vs+Bq�#�1��>2�u��r��>]ޠ���5�c6���Hӂ��]@��؊��O�0�=f��V��}�����^�kT���7�jdQ�� ��65���/*����p�5@�'W����Q�#��a��GpY�>�Q-GͲ���[�@����Uw������3�π�BJ}{�`���:=`D)�V���`#|��6jRl��qz��R��@��+,<�l�po��@�b��}�(���rE�ζ:�Wqy�$�d�tgHSZ�K.�B���A58�fl�F�X7E�:�g'k�b{�V��u��� (;�*�K�:�{X1a�ݻ��ʸk�)G��P7������ó��F����+������ձXa��R���ʣ`�&��;l����QO/��/��%q|D�J��3\����ٽ���lҦ4�im(qm� �F����6l'�g�U4����TË�*lA*E�U@![ڛ��N��#���8���:�E٣Q���+�]� �U+���La�&��c��ժ5��X�b��`�j�rș,Z�A��=���D\���ݽ��{��ݺn�֝p��g"H�q#�d6?X�p5��>�=V��������v�+Y4�U�����|�Q�B�"�`4ڜm�K5b�,}�T�[>6p�'Ϋ�>�p�_�nc/�V%JO��ctn���	�3)*�RNJ�M�g���ʿ1�
ZB=!���U�Ly����8��!A��X����vxMݘ�٢�&H7�*��U��G�4?�z�nɝw3��=���_��я���۠��ڙϡ���}��}��3�UN��
�Ul��M�e:���M����յtֲ�H'>'�#�^������2#��(�ړc��03T��(Cϥԑ�2[�f��:5���b����Lz��,~;x�/���cW�@`�#�﮶M)�b�VS V��u���j)�2T��w�>Y_$�CXg��r_i/8�-|� F���:�I������EC�-ߏ��a+�<Iy��D����,/��*!�xY��6�&SC@���s�$�N.���f~�jޕ-���ĆPt��QC�ُ-���_��aM��=�E���A�p-�4��s!	�,�;Bk�w��eTL�n;��fJN��[Y����S�A��;I��;�U˧�Wh4����E챛a��,�0���Q�����1˴��Y�;���EK��Q{1�q������ho�Vi����"�^��u���3���~�BK�86���s�K%4�����"���X����̴�k��pѥM���~�rj��B�U��u�T�C�d�_�)�=�(�
fzԵ�Z1Z��D��1�l�������.�0����VG:��B��y{y�Ƙ�:D�yIh�K��]��%�nϽ���l7&��e"}��\�L!SR��C�<_��Z��#�E|�����؞6L'��ݤ�Y��5��D�D��1V�m�޼���߈�e#�2���7	�;pI��B���}�E�-3�������N�=12D�3s�Bwg����&����0���4!��@�k�g~cE��Z��Vͺ���$`]�"�JT��Ǌ�6"�/��V����iQ�&iKXhSD(��-�O�:��M�i��7.�EvH([�h:���U@�����(�<�"��h�ѵ�@���~� #{݈�W6��V|�����0���}Zv��(��o�TEJ��2�7Xq�$_�������f� ��Fd5�p*�
h���**��2�͟�\07��N��G|0�H�>��gPB�I��H-����s��H������I:鱧*qv���������5�s��t����C1��c��x�a{"�Nגl\�=V�z��^�B�]����rJY-��I�R2�$i��P��d�dׯ9�\(��'{ô�^��na�DHb�bև�@��o��VبWCGY���u���m�ߎ�P�-�`��?�2.��|2�g�"Il�O� ��m������#�S�����pw+</]܇9ڿ���9e�{���R����)��T��p>�+3k�#�[
bVt5Z��ȠЯ���.�1k�v��}�bt--��!����j?1��["ģ���7� On�d�*�<���0rs�kjB\lL��V9�??f�U�E��0��h9* 	�,\.��^+NsCRr�!�2:�T�3�:����z��g��%��w�k5��	�������#O0*Vژ�)+k�6��N�=�0$Ҽn�ݚ�&��v	[Z�1�9��T4T<\��ǈC6Kƺ��jAߚ�ֆ"��K���x�)Bu{�Oo�1�}�%Osŵ�A�� ���#�X��L�E�7vi��IA®RŘ"����[sU��i:Z+�6�)��#��2%�[�g����ɔF��KY�ߜ�Q�}Xx4|F��~ ZӸ$>{����8pi��H+K��5�q���\�w���(��1{���ao{��Z��0���9�3N��@q�'�`�Q2Ǆ�=_gCB�(��i���\n�T�����h���!�J�	��A_*8y���G���۲�WEsZT��I�-�����,��P�+(�=y�lo�Q2^AI~�?�Ќ��ã���Ύ�h�H���1J��/wZ����:�,�:آ�aP���f~���G8�Z�[���Ǆ<�M����D���sS&��:�����]��F�����2Ԫ�?{�g�*��~c��J��~kxwnv��8xap�Xw� s�(��x��M�*���ʋ�v��'}�W#_��b&����A�,����[1T���3a]r<���!^Ͻ��:=�*����'\�/:�
���	&�$��.u�m�N��1��E�x^J�������Wy���B<��2����2 qNxy:~_�| |m��+��BU�4��1&3QL8z�3����j�(�R�V�#E�_�99(ʊs�k�{8z��dBrN��O�b��� C�"v�ܜÌ2<���b��&-�.��R���	��y�:E���U�F��P&�Ǝ�C�:�~haW�?�]�)��h��N�-�E"�4y��اUõAV#��Lp,�l��Y�d��7��R� ��R8ak�&��q"��K���O;#��&[���]N�R��?!V3���"��(q�L�"���q�0��g�4X�^�{U*���0T� ������L�9�k.`]�n]�v�(��鷃n�s�Y@� "zn؈dNyY�:Awhx��yWp�.iX�l ��D�9�"�N2{��pm�e.�͙�'9�q�L�^�M��ĀY�m��� O�W;7��D�ԺC��a���8�;�)�ޠ[p�fA��W��U~��N���_rc_�ĺ��v�w���g�!�/9�L�n���}&��YG���։��Rɣ����wv�Py����%�¾Ð�G�A^�D�z�����<��-������<{�E��� e�$�oӿS���$w+~��a�h��5'���%GVczY>$��	fTX��@�ĝK�H�diUͳӭ:�qp�k̿��(�.��f�2� ��ST�E����5���Gr>iRh}�E����h60�[#�:tԢ��݉�PA�M��?�K�Ї����3~c��w3N�m���@L���Y�2�t1��"���:{By��n:Ҋ��9J]�c/e4�u|6K�ԥ�I��X��;�:]B+HR�7L\DBQ�����M�&As'���E�t�d���J�!�| �������Py����7��e�;�h���:��7��s]"=@#�:yiE���W>���I�?`�@��r�N�_���qZK������VD��U�8�;�p�W��Lq|���l ]OL�I����ي�S�I�yq|�-��8D�K���A�7G�f��HOV&L��չ��	Z��C���fP].�>@DÒ�͏�|�]�Q�% �<� �i�(�P��g1N/����x�G2�`�3��٦�]�F��)���[����4��\���'���V��]��һ;� (�VP�:��ǓX����{�"�bV��S)�a�M>�E��L��6[eK��
]�=R��:�F̠��.�b��.%��-I��![�)d��};��Z�1#Y����j2�7����$�:������F�XD�����5�н�~0�OyG0M���H�-8�G ܎��g6�s�!�����J$�qL�t�TU/�g<XK�E���S^R��@*Ai��}T��6���BM֫:��Sw�Q������T�"��n��=,HB�%�L- �ʈ�~���#���yIx�to����=f~�{��&�k��^끗�=Y�o)�z�V��˪�*�B�Fu�� [_k� 2��{7S���"��ӭyȱp����mW^p=���bQ�1l%�������}ǭ��Z�[�N���-���$�{��0S�m"������Gt�O�{����o_��\{.J>�Y�6_�Jy� {��oԠ0��L�l���y�	S�$���w�x�Z�����E�i��u�$�ѷ���_�q�P�����H�JX&E����90�j(��d���pm4ͣ�ā/����H��:�斐$/���}ϻm>�]h	�D�ٚ�gM��P[�;�6�V*#����&ڂ�c틹3J�K�J?��r�����a�����4�
�d7Ó]0k�����+�����B�/S���'������6��e�������R@�*l��sx����HC�
s|I�5|^C��ϡ�Ĝyi�Ő�l�> :G���^��l�J� ���I,���^�zԆ���`�I�?͠�A�5q̬���	#����-Hf����Ұ/�Z��ʃS�YV�� m_�d���F��/��&�Rh9>�����q:����&� FiI��D�������Z?)J��j�� ���Е�5�]��>0��k�6�G�=����IYP�a��y�Ǆf�()����8���Z��մ���*��Er�a�k�/4��J%��20]j6��.�а�,���I�����	̽�ߊ
��&��I�18����-��;]s�ct־�{��U�)��Twᚗ�A˰�C6�wT!����0�n�zW�����;�Z	��A�T�tW=&dר� ��,�<o���*D�}�h�ğ�4Ǹ/���$�[�ql��z��GT	�8�`��|�k�VS{�J4���7OM4��{���B�:����A�1�JVac�o�h�-�U��h|��pv8"�hކ�gL��Q`��A�1���.d�!\�����y}Q���*w��ǥ�3wS�d�3�X
��&�T���X���66z�U�A( �dxg��,&K�*=W���_�`(�{Üu�_E�E�?&	�jJ��޾�Sl���p��{���4��+w n�{�؜�xj�y�Fs,4N�Pp���Y,Fd�e�(s2�d�>���d��F�'$9���
 ���l�d~U[_r-�,Ƶ�smx �u����N�D�BCz,����-(��R�C�h�CΣD�� �ƍgb�q���w�4��P����jx�jő|IQ�
�42�L1��E�����/��u���}��A�~uQ�~r��XE4D猇 ���2��& �F��h���6���g1?���fCñ��N�~wE�4s���������^��'���;}�?���i��3)�{���.D]�Z��iіs����/x[9q���$����-<Ī_�.�&O���A )3�7V
p�2��w�x�s`�Bʱ�+d�Q��˸`��\���&�L�R=�YB[�]�~��ra ڨ�I�.A�-������b�׼��q�s%Xp��)���h�U�d�~G~��� ɤ�:����Z��8@�&r3��^��k)aK|b�f���c���Q-,�S&,|�Qd~��W��=[9���4��s�kO-n���b���|�^�{Cm�FLc�^Vg��{�m+2���j�D8���/.S[ K��vQ�D�?�8�cF���=C�lM�6�D�6�T[J����ҙ��$�B\u'z��&��|r���ӻgODТ�'�1m����Y�h�Ί�M^�e��Ln�7v��h�H�̒4�v���?�[r���:��e��H��&V�����8p�W��HJ�2W�Y�7�-������Vڎ��ދ~������',%�9Û��	
,�o2���n(D9^�Ӆ��[����?Ҋ�\���� jͽ�<������a��D��[�+������$�%�C�.5-�����K�cȕ_B��v���hF������?���ز�!k����=o�( ^��&A�O,~+�O��ly.A&*�yC���u�P@�p�B�5�ݎ �G�E.4�����A�#� �m`�!��7a�2=�0@��c�}�bQ�y��n�|��%�5��;�=BT[�0����nD�VP��>�(p��{���܆�G�����;��>sH�.z�s�E�CQ���	ce���R�E�+Oaa�f�5��o �*�I���{��	}$5����+�p�ld0C
n��3�-k�`5�~��A���!1��a$?���8��_ �b����96y]�U����Z��Ji���N� ��*/�>��7�X�C�N��#����vU
s���aֲN�\�l�ox
�}5$�U�{�x�kB¶��^���@����e��&�
q�j�Չ>�-�<X��T�Y�6�Z�f'�B���ț��_Fꂄ�oj��(��F��%!Wr��,&'�宧|YCu�qE��v�A��p(sToDo���P���GA�$��C�)�O�CÊ�"��P�9��������yjۓ/�L�����K$�Rz0�<j^�Gs̀�F����s�!Yͽ|�0<O��i�h�&e|��k�����e�	�ё���i�]۹6�����rC�C@�י����*�
��ve_��'X����|��F7`����7��΅v��LB�?�+,�٘s��"�LT[+������E���iB�F��K�9�4��9o0]"���:��k��0�'��Շ�E�=W���2��>b��nH���:����DC��DqTSU���L�"�F��k@��rӧ�]�Ou:-e�a�v�)t�"�Ñ�g���ߛ5��9�M��"0H/�[��������ev�R*)X���éJ̦��f��j�{�E�k�k��*7��]dO�`j�xj��*�LM�h����i���`�C0DwI���,/ݗp��z��7 �N��(��?m-�uk�3��U��|��?�_�^��ڄ��/��zO#��I���ͦ7u�?-�h��_L%JGh�h����Z^�ƾ�ՓP<��[��6�K�0'S��c(���H�=q��c:�r���<��<!@�F�S)���ƙ���u��c:g,r%&��Vf�!��H��Ok���D�_d��w��ɢ�"�kH|�r� =�H{�F�]�w�1���M��V���LI���C+N��Ǡ>�c}`�sH���zU7T294ߜS,|���89X�~���`�Qn�7!ݐ?dִ�!�=$���_E�[0f��?r�0����b/��S�0�U�G�nB�������@��E�J�����M��C�����m��)��x1���k[�$�k��)e/[�N��et�2��W��!�T�.��{����P%���Ȝ����&�~Pq��Z����p�-���xX�Qu�5"��{�K�Eǀo������Hv�)"�Ǝ埩!�Б߂��@�'>O R�+4���%ڦ��g���t��\N�ݔ�i2�����U�� ӹŹ��
��EԻh���,y� ��(���{�f�k撵]�R`�q���$Ou%]S�������5�n
O�$Q���n�������������A�&�i�}�K_ՠ.����m����4-~�9xM/�4����7r�N�([*D�+(~���Ó���I}:��[=7�5'�;V���=ₕųuI�Q������U�C�hI��7�ȜK��-������~>��i ��f�5�I��	��j��cc�������y٣`�ŀ���K;A��}��^�a;0
'��e4kJ�%�k�K���ܥ;�t�)��y���xۯU�o��}�>E�K!~��V����
�����_-[E
�۬�nJ Y�}k�� �/H�����H�}�J��]D$PIf&����8�H�}F�i_��^��7&�Q�#_����j����n����QcdT���t+9HD���q�%���֣B�E�c^�$,�n�N�e��p�����w�1R=����ܦݵi	�e��7����fJ�JEF\���2C�{�%��C�7������^+���U7���i�����O�Q"��m�}�B(��`	���O~Vף��Z�8�Z0RlK�8a�ĵ;T� \��p��,M-g+|;e�PW�M�݅�&���J��D(���Bֆ�QQ�`�%��M��6��4��e��pn9d� ���흖~R�xE5�ч>�_Zo��,����ѽ;�ѕ���^i����Nf�z~r��)��b(g�|(���K�K�A��e9���Q^�a�*)��ˁb ��3�ݗ+���v�������>��2ҥ�I�6�bg7	��PS,��i͑����|�v?a�����6��M���&����7h����۰��Ԯ������:��@�aSx�J>p�A���SZ.k�b� �D�}�|pKj˱�?[&���C/J�|6�qY���&�ߵ��T�P���!�|R�iM�������K�o�����Cr�OV�q>[��K��V�=b�̵�qWZ���Z&̎|p}/�'���Pt!�3P۬X8qN3a]hΔ*�9%��=�ǂ��i�g��j���IҒ��b��¥��6BC8YI��fa&����ݩ���S���-֬�a��Z���5��bK�QPڣ^z���:�m�NU�D-"��8mQm����V�)���~.ml/5[���V�L!�=9�� ������h�q{Mlc��󞯳	���r�z�'L����e5=:;��L/b⎏���r�2������|��maǛ��Q,:���_��/,�Q�A+����J�2iu�1]<�a,�B$	��x���g1�z},@HA����8��É�.�v,+͵R��҆������CH��=H-P�S�*�X� ���K�:���$񳐸W'ƴ�k�uI7!�	�]�
I 9�����+E�8-������	9
��ъ��ǔ�u�o�R�{/<�;��ϑn`I�fh�s�2;�#��e�E#ӥT�
�;��]g�Y�<@��	Վ�e�����K������ŉ�T�5q��F-�Մ���Oc��te���;!%1�T�1'��4U?/�z^u��:j����}����+\�|�P�|淪�1T�)�	���9�KL�3�a�L ���@���q����Rc���&T[��<��{���^�a����-&}�W�d	���ݽu�DB��(T����r`v��;_���WO�z���ށ�0��xŇ'C�h��|�Fw^���U���µ����E|���f-/��(�	�U�崖W�;��XK#�{|N���`��h}���(;��+�=�i@��#殯M��̷�Pa�������s�w�����;�z�+��hY�u؞>I�l�,��S|U�V�uXr����I�����9���r�xW��\h��yRxҨQ��=	V �B�����F�u_5qA�@�ݘ��K82Xx ��?�H��/���goC��Փ�u��T�F��~O9 E���k�+�9�Fe0������ns�ﺰ.���8?���;�s�I��`�Cމ�~H^ j�.Z�"��r�7�u�>Q��U��Q�dlxn�K,˺��㏽/���`A�fc�z�7�G!�[��2��;�����u@f�P��Ыx��w����~5ߤ���R� lf����I3��+
��T6A������U!&B<>�w�]A>���^��T�h�A2�Fy����4;�vWҙ�%9m�Z|�߳�񮆝9
�{��UtD�oB
�Y��Uz�/t�8���<�ޡٱ���[VOy��H���(�!O^Eo,eJ��CRF�./������e���*o���}
ՙ���)Ȟ;�p��.���8^>���ڂ�ӈD�E����<:��"���1,H�nx#����X�tl�;:��*����0'@6Nf1(�j�����h�gz��V����a:tΙF"��<�H��@��i��JO��E�D�ϝ6����h}!���,�{� �3ŷ��T��9o9	�֙�G��!�͇L�g�'z�ȹbCt�P�}�B0ťgO�}���J�i�(^)��ǇC4C"�E"�dD���6�$�I��l	xzf�Jd��I�28�e�T\�Ò��fȠ����=�Ds~����)��L���f�J�k��.��.,ĵ�F[F�+����P=̰�&>��E�i9��c,�7��sS�߾�/eo3�e�o���_�۴�����}9�Б��ãL�-����Gc/'�g�2���8��g�ui--��"�=�ގ,tge/v���H�p�ʏl*{uM�qx�Rj���T��&j._�Qlt	F'�]+E22��x@�10} ��ym賌u/F����B���!&|�g5�V����̸�ټL�h�"�X�`��.�}���j'�=��?��=X
����!sq��B�bT��� ���t���XIm&x�D!]̍J�(g4g�b���0$���,���j�����esD$�vcL\>@,�\�z�jڋ:\�ӻQ�#qr�L;p�����|T��H�N�f@K�͢��?�} %��.C%
<��{	Ks�Dzt���Y�S�B�O���hx<7�
��]Y�c�2�Mۑ8���� �w�c���L�WA�OS��A�-kyC� �jڨ#c�����-�"j�-������hȝ>"Nl���<��}jj�.�(5<z���e�{�C��&%v���2����&s��Z	�X�݈�H�H����B���
��qbop�om�2F��3�� �K@B�S��d�?S��Ђ՜̓���a��$'�2��P��+-��ƈ��y�% _���@a�������ߪ�v�Ƹ�I��=��M�z�����&/��$+1��R�1I�K)�vI�C�&5��ƒ����n����L3�O5{��?��DmsfJ)�>���{*�g�((�KL� m	rc���`��\�h�������;D6�@�)p~�+ ���o�s�-��r�����$�?�4��`����c�������� j|�?T �mKTKe�D9��zάW*�(a�S	�q�~�����`����p���\��/�)b��AAgg�-�-_�Z����o~��`v-�8����
�$�ҫٹX����/�@�?
�B~�E@���I�\~�Q��Q��mB�Or@���Z�a)���"�|gL	�k�2����u�L� ���_Ȑ?��:֡ �ѹ��ެ!:L��A����Z�΀����	����O9�Ǥ7������@7��"3��K��`�M4��$�7R��tO�K�_1�M� ɣ�H/E����������@,�����S�SΊ	+�Q����]cz���Qɟ���uם����y�q�5v�!rO�qB3~�*B�i���=�N��eZpL��)f^�p�-j����P��`n} �[ɓ�غ�k1�)4��ebYg�����x����w�kr�"�&���?��! tGg��Y��UtM�����[�s}s��Q� QXd=�U����~��jnV��>,���ȃ�MI!��Fw&�~l�#�I�Av�J=�6{��$�}����c�+~�(��cn���b�6L�sľ�J���k����ōSs���R�ռf�f�v��;����-ǍHHXe/���.d���kûd�s��È�"�p�&���8��`î[6����w�0ٛ�}�V��}NX ���2�(�6a��3���	�nt�/{-���j��i4H�Y�*?2 *����`�����ֽ���c���dn_��n���i�+���Уa���!}�F��M��"�)��D�[P��o��]mO�I����Q�+ؙ-V=�_׊�<n� ��d����4V�op�$�����l�f^&���\s.t(���\q����t#�8Gz7���=w���IPJc�\~W� �TY8��-���X�f���m�C�����J�qY縿���&�8�k�n���b�����<�����yM�|ݠ��A����(/!I`ԟ��G��k�ES�Л1>wR,�2!*!�����0#�RcZ��*���wt�����o�(�P"�(�l7�e���y6��w�b��0�˃j(u�OM��RF&��WhH5��(�@U����:*pa��׀���]����wm:g�I�}�@�7�H;*DM�~�V�c��~�=�}�p^/z�(8e���a�֡w YxA4�bE�X���o/m�� ��:
�̛��zե<���V���Ǻ+�:��gDu�#V�d{�as�J���p/�k����O`k��+m�����V�Ir�G�O�ԇ;��O�A������~��q���ᒑ�n�exҒ n��/x\���R���a��}pJV���E:���?�k�$][h}2�׵Ħ��*c֡D�3W�/�8�-�z�Z����.
��g�Ec��J�O�X� ��$�b����J"d�����G�f�|���Le``���0�z�~��ܟߟ|�p��P���N�Hx���V�&�Ee�̽�(�vS�X+���
=�da�K~mN�t|�Tұz?w5�ˎ�z� �Vqt��=���^8w��7�}�E6������O��%�ˌ�cFͼE8l�̋*�7�����_T����`������6;��l-�K����·,��&o��7�������k�ةn�c�<Х������
J�~���'�5��5x8-=�%��A+��f��{�p�56��/qu��Y�c$r��+��G+�M��E��T �*�^��p)�Vw����r=G�2�@(�tG�N�oO���M}���m
��j-k� �\KZ��c����2':$����uW(�)8B���P�hw�N'�IQ���!�$������������2��������(�y����m�5t�����?�cҹ�>MY���L�U�K���K{�'ᵨ�8�O�Y@D�SyB9�N��?k5���
ǿ���O���a&�ߙ���pSw�:�u*G��a�쥙Ⴝ�U{^u���NˍB�E���X现���[DV���Q�9� �w���NS ���	⎔�MEt<��8��`c�O���K�˄_�6B�)/���W �� C��H�(=����V�� ��:�[0�E��b`_�H��)� L�n�LR̆S:���P �$���O��?�C�[��q�����qм��ܠ��V����Q����Cħ�p�*O�#�EP��q6�����0�ǌ+��N�����P4շo�,��}�E�0�p_?BfA�T�E�J�&g;\��:#y������^Y@@�_�9�"�ԧ���� �-���('����~�H�ӎ��.{,�!�V^i�B���	&5[゚�ɫ�7�X�B�ǐrdr:/������s�M��z���N��$�e�c�,W��뱰n�T /{/�Pف���{\���W�B�H��ݴ����2�����}*�\4U*��
��i�熀[�[6@0�?1-(=g��Z}��� f��1r��L���זG����(���C�V_��j�͇�ä��)� ����.U����E����F�[a�1[�a�>�F_�=U�@�#�_�M����<+�u�YdT�l��˧�QR�M���9<՞�ƨB��9+�>�7��p$pHhnc�#�������?��W�g�ݸf� �vҸM�2�%�;n��J_U��h��+m����)(H��}��en����s�;�Zg'��� @p�tB��^w��k��Z��q��~#��M���)ٰ�@���K��rCe�x��ٍ�����K��(�Q
0Ox[�>��,1O��it?���X%T�#m�ȱ���|���Fʨ֡cS巂����rJHnS���?��t�~����Z��w[�
3�2�l$�d����� �^l:����$�{?h��kW���IRn��p�ub�N/�\jں].�U$�q��Wm��2cTv����b��D������L����D��yAQũ��L䢯f���x�AummD+kx�J�fj\�X�Z��O���8�&^�)�D��^�Ӱ�4���?��9HϹ��r|�{����0��G��� �������|�
t�h�׈5|��>9	M׮�G-�4+�Tn�%�+�\}͠�r"_�O�rXe	Qn���w�=�(�)]���;��?���Ӷe��'��M%��䵁[[w�r���e�l�]Tm*6^�CWA�z0��8X��1��� |�T�O`�v�H�y�l��&�\Ӈr�s<����AE���Ǆ�� ����`,����#s��˪�ט>!L�ث�-��V�z^(�Ʈ\~��_����ړa?rV�;d�k0�!��b`�P!�Qi+��� ���/NI�ڣ�HO�Au�;M��%����кE��1*����9�G��,4c1,7�z`�����h�`un��6�8`��{D�P
#T��eɴF2�`�E�_��ePwչU=x�&��T�	�K�Ye�eGԹ�e����MȮJ�0U'ȶ��N�ᰘ�?�H���|����g+RA��QB����ʚ�<M>b!8��t��ְ�܂L�Nz2}���G���m���hf'��^I�Q�EA�~Ky��~5���$�=+F�OW�dU�!P�O�[�Ͼ���=���H���n�	탪`rx,R��$).z��.�?��� ���lb2�B���m�Y`6ț&i��b!"��F]JC������E��k��6q۪T����[8�c*z̥� ��wnM�����qٓ0i�9y��������~��5�+{z�EA�b1��t��`>�L��ef3U!�#4������V�^?�T�j_����m#	�y?��V�4U�E�%���Z�6�9` S�P�Z�(�w�-Ř�낏K���b�@��܇�[�nw~/��{��GJWt��K�����L��ź��ƶGJ�uR��=O&��o����P8�N�Є�sWc��=oVcoj��3�4EQ@�	���U� l��D��=��)huO�w�ϣ�
�nj*���i�T���p6�SS��ʽ�.0)��)ۿO�e�O���XB��rw?-0���Dy��ʔ��Ee�(�<�^?zd`��灠 ��:3F��1���䌷�`����x�~�h��R3���8og/�F�6@%/� 3���Bv.{p�F����;�t���U����*Ĳs!�ә�F�p.���HB~kи@9��m����d��n-宽+��l{,u��]�OWMx/�������a��o�6�����;�~`'[�G�*�z���im��d��0��:3e�_D=ܗ�I@-w-�O˪CI�	y�/G��F���tZ�P?�7v�Jŏ|��E�4�i�4�i��+���Ǫ�*�=�I�S����uyc��-S�w��RG��Orh(*ꢋ�B���K�������'�٬�X��O|-���Jt����䑳 �Ǝ �v{��*���w�N�վ�I�>Z1�Ik��V��Ƅ݌�Ǌ����@Z����W���,h�ɽ4��`e�ߥim�/�-ី,�%�����q��]W솂�G�צS�|��K��2���v�5(DP�Yc�I�����L�ճ�b6���vږ���I!�;�]����$���ݻk0�>0�Z�_����td
�1;�^T���{GE��V3?h�*�d�n�~�!"Sa��~�z��s�`,�!WC�;ZԆhUX��v�eBf�9Ƕ�����NW����_'�+f�3��{����<a�MǑK�*'2��"��F�X�]��	�0�(�"%� ��j��� V�.���V��^- �Ŗ�������'l����O6��.��Xl��L��Qu<XJ 75�k���`��8ɗ"洌�0�_�z}<O��k����Y��!�Y�W���$袀s�U��(�>�^ռ�O���E�6���t_��������/�	�������	
P\��Y��H��!bT��"�[(MA�g��L�'���O����!N[li�D�j�ߦ�֫5'ʛ�b�t��{1�����)X?#�K��^׌������C����Ī�~q���v" ��5�Z�Z���pqQ.1�a�7M褫�k�5������-b��9E��u�Bڇ���4U����zem�L�@f_m����'t��w9�Uؘ�L'���(�KOPm��I����bJ���T|J��c,ڇA�w"PΆH��w6�w��
G���}������7e��so��N�Aå���/�o��fj�`)���'&0����,7��<!����>�IÍ�p���w���d�Lw|���~�mC�/N�B	��9RI��Ce)��*�‘�{�6��A}f*�H�Sc�W�V"����s#�ŋ�:kxᚘ��n�_���v2��ް�AfЦ��1��O#C�O״�)�ߓ?$B�VH�<7��D���ϣ>V�a�$hsR<�0Y��ո?;P���z;FPo��{Bt�� �錇��1�]؝����g�GF$	�q�Q=��4��6y�St5⬲�ˍ�\:Q��?Ul.�sc�(���{I$����������eM���/X'��'���D�f���w�	Mf�����R�x���A��}4�1h[F���Ե�� $�t�	�p�4�\ɤ���«_zfs,��OK�,T�����Jp-�_<?���3��0;&�K8�+���01X�,��'��	�E�LΊxU����)�I�P��\�L��I��������%�QNP���h��4t�r��]�k�N�v|@;�uar><�����I�<}�[�Llࣧ��ܰ�":�cUj�>y)�m�J�x~dI���j8��`��
-�d�� �ђ�N�љ*��c�Y}p&3�����S�N��ܲqS���m���$��� �yr���6��|�ڼ
ҳ���J�*��ć;���xƶ�]O�sT]��Mݐu�!\��D۔nd�N�>�B��li޺][��P���|4a����yky�A�������S?9��\����M`f	d9����-0�?���Ow;�]� K\�xw�a�aV��T�5�d�g��n13�'C�Q4�R��c a��G.�cdD!�$V�uA�}��h�&Y��:���9Y�xvSs�	�7��(�	�^`�/#�Ȫ�P�����SB�� +���9���\����dM�����1����y�5"�Z��n��#��d����&i�eu����$���5�4�`��I؁A˨Q��=������gR!Kl�k��W)I9�����**�Ldu�� 	�\72���8�O��݅P�R�*̼$����7�|iv�[s�njW�H%�d�=Wa<���bx���#B*��l%p�lgV��/���~�U����i;�j,��x'��(�8ޡ�%sq�uE!�߅N�:�z�`�7��f�$h���بp���JI`���=�s� ��2~���~�)��/U!T���k�(�<,h0�B��$��f^H?TOT�-�6�*�hcOq�Ā�Ɍ�O*�,����^�d���/����	�R)Og��F�C��Ԧ�psI����L������뵚�+0��s�U�S3�}��9#�a#�m��p�-m���>�d_q70<q��3�P���N���;Eā�!b�m��"B��?o�ՙ���J��.�T�����	q�_5�[�X�i��,����Xv��y�H,_F���X�����[����4����܊�l�r���쬓
�׀�J�d!w�,ۤ�2�gt\�2�������*� 7����5��E+pSݾIx��t��&�"���(�5�`��_�<�%o�"#�X���l�{�X�i.6�c�~����BЖ�š�W�<xD�`!}gy���v�/�J&t�,</a�d�".)4_����5��9��0F0����i�ư���e���P��Rc�� ~�.��IZ*m�|1l}���S���F���Ds
p�uy�T�;�O#hh�=�����S� >.ת; �k�z�\'S_����d�*,�Gi���?�Pḍ�d5����#>�g7>7�](`�^���\Z#�B��G԰����n��.����@'��6��ŧ ��0 �����ȅ�-���X�� 
��V��Չ@$��L��r5�,���I�r�K{�9�vj�GC�m@JKt"�E;	����%}x�͘'p�a{����ɦ��m�ׂ���JSr�рﵡ�L�o�_h��d?]���O�Q�rB!���M]�n��>/�� ��:l�9N)��w}]a��k<����%�U�Ⱦ�u�xj&�s�|_6U�>h�����I�[����WV����$��u��(؋��7^_R{|8�~�f�䘢IG��-�櫾x� r=tU���U��f-Z�K�^�p��Hi�ao\��BP�����B�����G�����/KS�Ɔc=��]�'�%I#�H_DHĎ�8����gQ��Q
�q*t����O��Cg�Rqķ&זs��0�?��|�"j#,H�~E����k���#-�}%}K}�#o����~�$cc1��[V8��A�P�gåR��ې/��mh�Yq������sH0�0�횼�<$(��g�Wȇ����~vH�(/5b�ZG�Tg����dF�#�RՒp��2�R����i���Z�}��_4�W��C��|k1�f2��ta��[c���A��A
�4&�}������V�]wv��haܙ?�f��<@Ҏ,�Q�4P�۝�N
�`9���~pId�/��
�&1q<��4gFf���ku�=�!�:��i�\DB��m;I/�ν2�ilRb�s"ia�f[<����5!r��~��q�ݘ��s�|	��'H}�N6՟��
����W;Z��u��Pf�n�rF��Go���")ܕ{��y�y-�a����4�k+<<V?�>�_��݉�r4>Bc����t��K�t��)#�E]��Ӄ�Rw������״���s�9��& ܼ��# ;�Xg�ڃ�cQ)܃�ݐT�\���a$�V�qûK�Zl��x	����]ciX8A�B �:�p�/��EV��~��bo�4YxD�m62�a(�S b�>d���{	aLf�<�+/82}��0p+-~րkb&2�U/���;R8�}]�Xv����ԑHaF��]��>��K���X`���9�Z� ����9/��U�m�"��pM�*̿�Oq���u,�O^�Z8�4�G����n#�H��/���@�R���W��S�&a���ބI�U���ݢA��WuΒJF��UM��n����qڗb����j[7K�(�!� ����h����&:5��
[���2V���4�Y��1q�}��e�4��G�uZt)����	�VC������U��!�p���02 �k�|�Wk �Ӕ�y7~I�kU�!�m��z�QO�ĜH���X�&3ED���5�V��c���t�U��IjN�sl��!ԏI���`8�;�v�I�`�)��^�F ϓ�h��t�_�n�:��'jz��^pR�x %�T�Y�kWC�����7��c?%��cC���F+�[x�C�+ˏxWqXtr�����/^��&�(N�J��c�-�u�
U��{fe�#oh�s��ԇ�~?�b:{t�1�{��_y# g���EㄥRĲr�>x�I�6%��^�35�u�Xa��ԇ�߬<��������2�b ֺʎ;�6�Pt$�V�Q&4�h>��R�� ܼ]�w�ʱ�����S�RX3b��;r~�y�5�u��}��
�2�tb���;^.�Y�I~���ۨЇ�祥Q�O;�����u�����1��Ӻ�m��J�X�؀��p�:-5"���ۋ��1&H�,��
�A��.A�ɽ�c�!���9��):����rm&�?'M�H[���|�#+�$1�s!p�fU��Lp��6�H_�$�-�g ��΍0+,ǍYW9��|tY�?I��֮_*������ �9[�o�9;GV�<,S�'���� �u`�
�^�������Z6	�:1o��a�"�q�$~b�}S�?�xHn;�qJf�~�i8�{��:KM� B����M*�J���p����;��XJ�S�'r��#Q�����\1tbp����O[���x�١�P�A$B{;?�^�g��yV@%�#���hS�RoԮO�D/��K�#�)��A������8b�^���sv�T�m�()T׏:�Uc�i�=��Q0|X&��Y�D���A���׵�փ�4b*&������ތ�P�n���q(��c�cA���y�'˹�7���u���w��o�؉�'���fਔ�������V5�>>�ڞ���?�?�;�{W\���s��2��1R΍�Y���{�M�c%H�U�\����y�ru�2��S%��Q�weh��[�	X�SZhc��mƁ���7t( m���!������1�'�44m\�m`Ȉ�Psf�Sl�Ԫ��'V��G�򼞲1��������Y�4�)�w��'�B�o�kc~:���/�Po�#̍�L&w�4|��G�-�U�a�tZ	|�b�Ml~|��� �f�Z��%�����<U�q#���'d���H���_�Ww�T�h�(�و;�6���c�o���3�f*�\��s_ղxi"���xթ?�BЕ测�i�ڈ,���u=U�S�,� ]�.xhI�#�)t��V`�Vt��-�]�����T�чS�f���Z�;^2��Q�$GQ�wWh��b���d�Es���b<�]�
	"D��xd�g �3�[�ϣ��z�FO��1���\mГ I���	q�XV����>mCL�9 �T�:�f� �s��K�ןؐ����ӑ���/�b|�)�9�|8Sd*l��+y�-,6�-�u�^�!@�&nI2�q�b�ߞ(Qg�t�=q	��l��"�k�z��@EUaTT�����S��Ė�� �.$��*�ޚ�I6�Aˡ��ɹ���͟���$7BkT�E��N�)�xQ��W=y���!�;b�>�l��K �ڜWW�GX�FA�4�j�Դ�� $�-��F���;��s�Wo͛�8 �4��d�X�{,Q�7�,�i�*@��7gPȧ����<X%��i:z�>|�N�|�D$��+-�~��a@�3E��R���\�WU6���:�j�/��iȌg�Q�	,�v�|�w����o���*��������1{����oTu�#~T�*Q8�?��'�?�B���aF���ͦjՆ�k��wkB�)o54������r�G��c(��M&�mB�mn
�W���-�_��D"}��`��"�WK̵��<c�'� �禂ѱ��p�A�9(�v�������]��u2�����ѽ���)oC�Í�)�3!g^rB��F(�^�q=�3ؽXO�J��A]��&�X0�Ҳ����fR�^�~��f)�l$>�wNs�܄$ٔ/]V��*
٤�@�#�A�H�!`�g�*����z�ގ�/�ۧ�`�)���3��'c\�G��Xq��ut:I�Q��c�C߼��)���D� 2 ���u����V-��&6��˄z(�r{;'Sj�)�����8�^�>�:��P�NLG�H�z܅^�ѩ=����4�u�vw��tq��ɩ�sH��<��Z}�����=�hY��s��ѕ�Kʋ9�L�b~�����&f��^�_0i�~+"����g{J��C����]뢞g�D���<�͆^�ʫ$��XV8��AyG�-qH��hl�@���MU��{��-r�/�e�x&���1g��M�HD���tAj��ϻ�5yl��6�aBo��u�D{��� �=3��9�����i�i�ɯ�_�f]���Q�y�Fb�K�Fg7�^���wb�J�)_�FSȷ뺴X{��%���GQ�O��3�+\D`M!F��N��z�oE��|'���ӷۤ;���^#G�����M���.2z�P8l�>����1K@*r��(�g(�]���7��-L�W��+I�.��M�S�u��<�}�t�l.c*��c�P��໗�2��C��)��~�gF���{t�i#���92'�dC
P���fe� � ��]�� +�=l�"' 1T x��8�����`3��aY!:-��ơ����z��kFG����V�"s:#CW��k�Ԥ�s�M>(h���.s:�i��q�˺���p!�Q������k��8x`��_ۦNg��0o֖��#s6������e�>U�4�Z�k��MT����s��Ln�Rt{]C�7��ؤ�P�1������Ԑ�3���+4$[��e���@*(�R���:e�'l�^Lݢ�#Ҹ���>��mm4|�T.4��OL]D04u�c
��ɟ:��Wϼ̌Z�-�ې���]!pd-�U4�NA��w�At�=�k!#xVȣ[ӀY{���1e���@?�H�s��	��x���g���	�8>���#8B���(�D��k�Q5#��t�n�<���M<4�����~G�r�:�. �K���,�w�¼�:d"KPW�p6a�q��_��������*c�U=PnUB�W����M�|B�Y�)��A����i�B�K���� F���z^�� _�M���܈|(&���Z��"V�	8w[����4}^h�.���kcY1+y����ro3�u�i�p��:���U?ӬPߡ!;��F#�k$s�i�p��1Dc1�$���NTr*��e�z�-89�y�9��:��3�S�L+�#M�u�{��5u
1���xe���K����G_7�����u����&!��G�}��(�s-\���F�� )����W�$�Z�]ޥ%"�$����Z��{��X��� �q�IN�ք6!΋ހ�ƥJ7؛0�![Œ��|?K��ė(Pn
83�i>0T���s`�'�ۆ,|�'FD����:����lVP��?Y r�B�m��O���>מ������a��v�����ĝ���ڑ'E�[3OR~qZ3�7�.�MK������|_5��{���%D�����|Nt�m0rC&��~����Xס3�~�~�`�EvZ�eΣ�#=��ɍ5���Z����L˓m�yH��li5�s�A+`1�~,�f�b�T�V �d��MT�:��W��{�N"�����L�R�xtgo���E��>�g�)#7C����<Ą��l�@ ��r��q*8?&�Y�ӑW_��0�t/�����H��U�l
��-fd��V�z���?>�S����
(�r�1���� ��ZW�u����Y�m���n>Cc\2bT�=����G��diDY�.�>�7A���9gb:��=7��!'�o< �KY%�8�2g;s��y�yz���ZI�b����#�����q�F6_����g�@
#)i��XM����Ivo�l+T,��(db�E��H�!��y5�R=SEӱ��1���t�l��6��!C)|A�QYX�2�ǆ�� .��"��pJ���,E��*5isp`�ЅY��4��{t������5�� ���T�����dOڮ'g�'��$h��3?U�Yd��Eo����%�}c2{���!��A�&�7�}QeW4�'L�u��G
4�ϩ����n�������L�%�9��#:8�˖}	&]ٴ���e�9����	ZKA��n����
��z����'Tv$Dol.x:�B+	pTy³TC�[¯�eN	�cA�QWh�y����P���Cn���yJ�������솟C1�+�1�x��²��� 4�`��j��.��"��[e�'��0����7l6�~k�qB.r��"*3켒�Rӗ��fް���Wπ^��
�b�����4��� ���I^W��w�&��u.2Oe��ݡ���/]�VX��~\��AU���R3�c(w���k4��o�.�����*�4dM������l!n7�G<����3u��s����[�~	ߩ
���ا�ߢiU��p�V#�C[ ��m�
����g"~�O�PS���O�%���6�W<�A��IB
�?��b�Pw}b��NFj*�I����'�U޺P��o���$mV~�e�}������0�H�7c�K�R���t����G����8M�� �R�Zy���Mp􌙝K�z�4�]�CT��fV1��,DT��f�v�F������"��c��GJAj�m�4(Չح̛�g����t��KHz��I,R+�@E�ڑ���G�> �� w#�:��'3���+�7?��hot�<�F�+w��>�2��޴�oTy�HR� R�Ό��p�H:U��=��?�0;moE¸ #v�7��V�8��	�:KPg�Zܱm R�B^��,4y��6&�4�j@0Jj���E�e�(���B�n`���*����1ϊ��� H��B���0�:!�#�71G�R{,�~��͓����y�؈I��� �Bꝁ�}�)�'{�B|t�,�c[V���޶��T%�%HQ	��W�2�<?���?���	�s�׭r ��q(�M������o��/F�9�D��J�������r*�H��=咏��X�a��|y�Dy��z�҃�z�<��i��3\B�#�@�;�sϏ�#��H�~�m4� ���wjRg��$�7x����`�5��k��6,)�K$��;�Hv ���%�`a���F{�����؝�{��?��K-��~˩}�l�τ@P^W��Z���0�s5�.#2������v�Y9Ui `��������ה\�g��[�0x�	�ҳ��ϷL�� ��wm6�[���hhvĺ]���z����_��~���g$����!���@2P��T�&��b;�^3YZ-�'�Ț旚���$����ܔYo~�����������F`f�u�b��o!0p�^��!6�v6Yn����lAa���?Kz�*I��l���%��KW�����^��ADb��?5��uP{�ku��&[9��Ƿ1 �(����"�Q|�
,�|f�|��z��!)�{n"e$��Ϡ���K����Lz�3�����ߑ�2Y����w�Î��G)�~�GX��]�dL�9����O��s��(��{�4Sv�C����Ʃ@O�N`�	�O��픏8\]Sf�zV�(�P���n��ze�|)Fq����pQv�l��X5]��y5�"����vl��*��k���o #�v��K>0~y\�x��O+\��	���>�2��7L���wڦZ��+������kEn)
u�H?�xˑ���F���kg�k��bPY
�Yl�m\R��@K_	.w�7+����RG�ԓ��� �S���Xi����W�}��}-��"�����R�q���C5络}rP*;�l�����n2��nL�d�!
���d��9|���I ��74?-�N���[N�V����*C��q���֍��˥�$(� U�1���UdF��y�W�3�y�=��N� "'�Lk~n�.u�#�q�U�9��M��k���ιn;���Ğ�V'yBF4���vp�����
v���@�[�a�A��n� ̆�	Ϲ�o���hG���:����M �<�YYZ��ظ�]$x)�!>8wY�d~ �N�w^��/ pdT3!��&�
���PL�����H�&�_q�0���W��?s�ܧ�Xwjd�D���D�=ӟP��u�H�-�j�;�4��rM)
��BP6��󬵻��x	�����m�̑>�BQv��xJ��xO��1�ʮ���G�.v�[��Oj�q��"�9�rq��9���a��4�I��)��ϔ� ��b���_I��RKR��a��6�ҹ�tŇU������\I�ܸ�P]�D���)#^Q�Yg�@}QHw��u�R SJD�p��@�������1�c�+��@��!Ɔo����z�����h�W�nMš2r��a�r��j�� ���A`�܂�7�̩l
�Q'���Я8G��\X��-%Jnr(��a?MF˷o���ev�O\�E9���ie��q2^�"���+*��5�J$�R�}Վ�3f����w��D�et쮺�I��W�C��P�Q��z3����1��HA~�8�ڻ�7����߼s�}%bE?8~�3^^��E���7w�k7%�K	곽�����@�t��h6����1B��Y�~���#KMv�A�]T0.����Z^ �9= >��Tϫ����ߙm�}����^��M�0f����</Dy�4�7���Jm��SXz}��Oq\ {%�gK!�GY'�@K����X�k���=bE;�ėC�&9j��t=S����,��cP���@Y\Pe�`��r����11�b
k�G�u���(��M"��oiMb9��� X�`7a^��gD���O�h
0��:$^"�au}{��UÌm��>TS��-�)�@7���-e���)�h���W�/
�k%�SPg����x#cP��ݵ5<B����&#�*ߦGf� �$S2u!xu�z@�y�� T�5�3+?�~��:�[t����b� �T��}�?���bLt&m�\@����#.~eJ ��i���,�Z�*�W{��gҢ�m�I�Q��޼nu!�	#Σ��2����oj�������vnk�+g�=��g��ly�)�27d:#&��?ͫB!��@�(�v{ܣ�����N*��ak;��_���/L�"nf�#�mt<^�䶢����r~5�"����{W<o2��>d*�f�7^*dL����ql0�$��(6ٯȗw�#�n%%Uڷ��;i�F`��0!+ɚ���X�?D����� �����	�s+X��8釬�����ˮJ"�T�wIi-nҘy]�E��^s��U�%ȸ�s!P ���`�ZS'��'Th��v�&�6���%E�u�v����{���׻�p��6��K=t�HB㸻��j��R.0������[%߸<�V�*A����Lo��4J��Sy�
H\5���{�_���Fݕ�S��H���0r��,'z�2���p���U$��u"yH�V�v@c�ԥ�u2�ɏ8�D�0��P��z{ZoځF��K�rN�5�Ƌ�_�f?F.�(��X�;����^�%d�X��=u���h8OW�5sv��7�mڶb���ר^�O��O�Y+���O�>��ݠ��PS�(7/8���[�	�0V6Ԕ����ci�|����{�֜�w�& �xP���Q�b�d�k���JO�,a9ض�Wp;nB�%dk�֐(��n�(}������F^��&6�7gۓۏ�O4GS�a��iD�'��%����CA'��E�(D�
&�m}c�ox���Mvd+��ʧ6�_��@�"�ĸ%� Lo5`做䚗��^�0]��E(3��)e��<�ɟz��C��5y9��:�ٿE��Z�mv�&�,�pLX��:�ex���3�O�SX�q�{�1��ѓD\À�";W�fQCR֊��fe������x���`�:�bwDu���d"����׭Q���g�BnѴ��7�����u�������Ǻ��>�pQ%�ӗSwD������Ywm��V�F=�� �5g�ͨ�'����J>{p�����¬�X��W��B��eW�*sRv~��\�O��NEm�@�ŵ���2��@���������|�)��J d#]`�'�˔,��кǈu�~4��W���O��m5�=�nh�+�n6S��C�ߦT��d�X�IY�B8����ҭ�T���J��m1�d�%��υ��X�_�w e��c�^�(C��߸콳����`�׊�"�W���4#��e4`�����4�l��TA�f��uU��7�z�|򊮥\��]0�7L�
Yw��(�r=zCZ.�h��Ϭ&�������@l:�`*�J�EkB?��]�R��ӰI:�>�,c>B�w��O�qh|�U��p��IvV�0�`��f^���^XS`���E܌��'R�~��(�A sL�A����{o~��p鱣�I�q���kX�����
KX���W�RK����v����)�&G�)�Z��q��{T��E��ލ'��#)���=�"PP�j��	~���]fΓE[�@"K�{؛TJj�������:��#j�H��M��޸}y�O��O4�I�J��6�
G��I��4�=��7�c�Ix�R�[���N�(�U
�<I���څF�կʫ�ԯI� �9}��-&��RU��f�}1�*G��"�S��ݟ%#c�	l��̫��I8Sn���;L���r��y)��XQa����_4����?�]�Z�ÿ�2>^�D��dvU~n[5)�_�|���=�u�G�~n����X_��}��bx�tG�P�����H�<N'MvlQ]���-���,q�+��q��|�D*̈́p�W�r��e�������z��g���|�r����@^��m�o�U ׫Nie��M ��_����Z����=������)Ǳ������y�5}9[�5J�7C�9�?B��I5Ա�UJ@aF�N)h��,�xy�ߠFd��B�����+�L	d��P��d{��
M�8�2�>Go�
��k���,g�XN�L�tR�sB��3�ĝ��i�hc� �q�9�/������
ͭ ]��wA���8�)�j��9�e�{���f?�~�%Z�~�� �:��nV8-�S��N��o	�Mf�f������)a�>-Z.���_N��_�HX)��M�z�N�2$��$���0BS��ت�{E�t/����̨^>�"eiܤ%���8��%�*_���Hok���r+k��
��[�}��L�~��K�=0��'�*���?��Lx�ظ jdQ����A�zNA�EUٓ>�l(����V�n��KS�&K�`"��1����U�\�6�{�s��Q�8�Gu�z����� 
JTf�uv�_<k�P�_
m�ZNt�0!1�Fu����YL�'�s��m|	���Ҽ��?���`�)R~puZs�3�v��4Һ��@���w9z�_�~ȱҌ޸u��h�w:|ԗ��O���d&���4@iM ��1�N�0x�=�Ot������,=�>��jf�P�ɇ$ �-�/����B"6��n{�C�3n��t�������2�I7�/m�!yӾ�#�3��j�|e�͇ bd��$�+)������t���Ѱ��m�iA>���6Ҿ���x��;�YvZ�Q��a
�U~l3%��>�P!�0��ԣ�
gm���Zv�p'j�W�Ҥ@ĥ�0ׄ���?�g�	wA��a���m"d�G}�T4�4ާ4'�A��n�(�tR�&��F'F*z#�����u0�GP,�r,�8_���WM�(ƺ�Qpe�7Xx�q�<��NzN��/��=�>�h���y�?�WTk����%��H)H���������H �q\I�xh-U� �6qA�Y_q�����;8�S�ߗ�ӣs��l�|J�T������ЩB���$X��j1�kM��ܫ'��y�mAP�x�����c7+	P��J���C����8�T�5��H��{?l������9�5=�!�D����+�z3�g�Jg�R�$ebO�hқaTϐ���F V!�������Ye�k����.���`�K�����v�����łit�c[UK���`���'*�CR�E�� ��̹g��2=��nog�~V��Z'�u
�	���]~ܣ�����{�^ѕ+@��א�o��]6i���	!Ñ�28��s���tldnX� ����#�����گU�����
�O��o�&����$�����%�d��z�ߔ�>�}��� �����&����{Ρ�
�"l�P��]}����R_�<�Ă��!w@�k"xӛ��c��)��U�ņt����XX+����H��
�"��ev�d�o䞚C�L�Y��׸o�ũpq����D����o�����A���
��/�w�֐�>o��OQ�̖���l���Tn� �y�(s�� xM�>N$��o�+`$�0�����Fyk�d#��ccߡ��g��Um�Z�n�5�_[��<dID��h�۵��HkIj�
^��q��y�Jo�Cz �F�T"ɘ�$��z�������(1��XgCL�g%:0g����ν�qil(��+G}lf����oF֖�h��z�N�� r`5M@Q�+��d��8�+,��� ���9�ǧ��sXv��ר���B������V�u���x�8Gw�V֨�+o;���_`Ϛ	8�7H��-��QlN�t���h��k	�} ���n18�!eU�}��T��ZV���q����(`�yZ!F��Ϳz���Ŷ1r;R�B+��F�K�Wp\�`�Ī��[�*a����t�6Hл
�YV�� �d�rw�|_?��^*Fa#qN0s~�`��x�/4�ndX|�P�=3�۞ѕG\u��>��~%/!,cA�Ժ�55lT+����I�KO�j�s L�ɺ�	,s�kR�'D���+�������V��|�� �w��1�tw\�RJ��z.�&2 ����&հ) M����9�9�D�Y�ṇ����zhx�V�*H�t�||�_��Wc��O�߳ �`J}q_��cJ�������O�t��T�:椭�#� �}���ҥ��"������7�ch=���`N_�AH�05#�Nφ`�F�x����?��L�E�a����Ȍ�����Mz	)�ΩV�SdC:��?.0�;m�i]��3���s���Q������6�|�?Fz�@@�!(#(�ߊ%Ե>:V�]���U6n&��@�eJB�i�����L��Tuc,T���?.l4���(1�NL�$n�d�őG��c���6�"�
QXJc�@�騾\�[��� �@��L��<C�.y�epX����FsewE�숻�iJT��A�������jR�_��gҙ�(CoŬRz�Po��=�#��46>�0+���kR&s�&��f�_���2���3�������|�`�r��]��`�_1�~޸��ؚ���m�8�dH�R�Z��	͓x��*�y�v�I�0=��F�	>S�E���#�97yy1�xj5<�Ṓ��BbÅ,`&��D�a*����~+�_�ޤ5��2��֊+��IB�U���f�� �"R�|'��}�����K��*[ud��\L���صȺ�)�C:�5]
�U�p��M���Єn�=����hK,���g� �!�{�|;��;����=776��)��	 �;f� /����j�zTU��3)U����{ùo��sS�(��"B'z���y�m��Yሯ��%̥6f�s��t^U¨�?RhcH�ԧ4��xg[�!y���2��&��#B����9��ː�"=�������kޠ��KQ?R.�30�j�x\s����C>�֠�l�8
g��
*9v�pI��a������K�q)����(
҄~l���m'唕@=���yݛ�+@���u��kjN?�:2H�3k�'�����W����(kM���${^q�x�γ#�L�"si2�p�W½>E*�XD� $4�\f&I���5���_�˃��,+9vd}{.��\.�U�r1�z�d2}����կ���2���)G*��9�ʵ$�%�F����Z������Kf�#Q7�}/%���A�N�	d�.��H��G#pOB�5�]8�q��+<�JD�XWî����t���{ȉ*swmu��o������j���V��'�(��R�*˛]�<�9��Y�R����n�Rۦ#��t܍��ι4	�tG_�/5BR"�
1{#D�s�wVs*�b\�=Ƙ�o��yF��o+N���.�$�MO�s�v��<��|d8��)
צ.̮Ȼ�g(T$a�).�	�M��Xk0Se�t&�e��W�%-����y�)�EA i��Y����-��쯕dlH`ZX�_@��-��Tl/�D��q�ܙ1#(Y:	qS�7E|T7 �o}�U~��d��my�$�b��Rn��k�x�"ڧ��~a����P#�杔�8�;�OkPb���7��;��-!�U2O��������"�;Ms.U�a���%r�>Yj^��HeV��ߖ�vOYh��Ǔ��㩊E��A���kP\����X�F�^�w k]7�����fF�uT�k�UT������T�X�Q�u�jA�7�?2y{n1m�Mߛ�|}M��;�x���8�H������-f��Q��Z,S=I�ms�'G~R�֓���n%��r��� ެ�Sgӵd�6�3��E�#��C��:���;����v��}�C�k'��H�/��bY��>��nx��o���֑0�6�� ���>��5�٘M�X�ֈ�6BذO�H.�NP8.�o1`����@��~[�ˤn�X��eK��\�oKQ��^�����D��0FD%�?�Q�͕!���x�;:�$ڼ<"I�<�ǌ�W[X�RR�0%���������k���4faG���������!҈-1�D=f�����\yx\Rv��m|����6:����X��$?��C�07g����J����N��x����/5(.��p�i}���{.lZ}�0� ��R~6�Df*u5�����`{��vιR랖E*4=�{b^+�e���bH���C��}!���,����Ĺ�}�uol{�ٍ��r"J��1��0?0�Q��`�]�V
��-�==������0���E66���B�g���n�{����zbڰsP���L��?d!��M�5T�{�
�6�X��bw��v���mJn4X���[R��p*�D>�����6�ď���D5�)a\Ò�����GE!{�^�O.%ỡ����e��6�plʫ0-���Ҥ�Nŧ�̆�.��6���9n��-��/��#9�W���[��j���-����V�����|A��7��b��v�h��Wo��Ћ�t�xPWО�!����&\S;�����YQ�`��9�W`���,&�▞k�H]��5�u����J
�d�=�QIwPu��M@;���E��P���#W:�F�q>�j2 ��ʥ��;�	���i�W������La�YIey�����ǡ��E��&P�"�Z䡤2��(����(&g<
+G�������xց��O��7?�T Oޣ��b�F�-����z������H��� g1=Ժ���mS,aF�J� �0~U��m�M����=���r���u�bRe`y��8Gl$U"�P��4�S�6��L$yi��{NP�5�N��1Y3�_����5�L;��׳�NUFj�m��Y�
CwPFйס�L骄 
q�Y�:hf�����e���SL�&u1l��N4{\��{׸��9�+m8��}3�s�B|�F�J����������|^��_��I�{��������������n�oD�׀c>9���Ǌ<3��|L���~-j�X����v��͵����~m{ͮA�+t �����A��pg�1V7U�.�j��|��!;e�-�s����}�H��c�˿��P�G{���|��2�1����B�����2��`c����*���-�r�m�lRk�o����ś^��KJ0^"�&P8:t�f9���9|��%I"�܏���W��?�62��S�i��*��ʣ���S�j}� �N�=
��J~B��)��%�$�Jq�����EO��R���N6��˞�ww�:H��r�Pp<fh����r�B����am���K�VK�޶7�IU1�I��T+�H�Du�e�(�-�Z�\)طF��^+�����9Ee�	l� ֜��kd�+Z����W�i���>D��n�,7�)��ܩ���W5�:s_7w�Q�<���`�9#S%�M�=&���{���}�g�P�Ǵ���@s�����t׃���<��:-�k�H���R��%)Y�rE��d$WoØWsb�{���� GeBG����-%9_������͍�$(���T&�C ���eum��|0�#�4�	��C\=r{�m%�o�X�Oo��>�- ��W�qiL��#��,۳:s_B٢��Z�f��
&4W�⥮쑾����ݙ`��/-�3���6
%2=U!�p/��в�٘��DU���[]=�9�e��m�>A����B�s/3�>ۗD���c�&�$���wqUh��#�Ƙ�I��!-Y6d�E�Hz�OϿ�P�{�x۸�!�P錆��Q�ЄO�F&	���W7Z�BcD�R�d�������n�%}�"P|ff5����Z�גvMR���.�������U�|��^���y�qH�Qߣ�aL�Rl�b�+�)K��YG�Z;��nl��j!}��8�EL�i6����������$�[I�>��:����̪��k5���vT�$Bh4YN���ws�,<�@;�<�h=�PZC2C����L��2�	o�8����a|:�б�z݅�/Y<K�M�"-��R޷�ܽkRNWܦ� y�ҧa�v�	��H�5X���I|3#�,?��ɂ˒�������
	���lp���G�S�9̍�䩲~�+����86�/E�/}��Ҫ-q �`Kj	^'�~��!����P)'n�0��l�).�᠅{6v%/,{���"��a�5ٺ�B%ׁR�X1�T���p|dHvC��9{�<�=d*v��OZ�5R���=Z�U��w�3cZH��d׫�PLÏ�rھ#�[�.�0�{�,�$hf�GՊf,ޔ�[nl2������]��S�Е"Y6����Go­9-���3@;	Q�$��M!�ۛ�Y��S����<�=	�rE�����AX ���\}V�@����B}�~D�-;1�hdV��QP�F��n\×���_���sx������b	��]�ʍ����[-8��K��,H��,���p-,��4/a���Ie'���dl��e����Yh�U�]���٩��`�*�Ia���b�z�0]h�a�����N<��ܰf`��}N|c�4n%����n]$P$;3
׹z5~�$��5��W(V=�0�'��U�G\�-pQ���4V�f����� �ha;V.��L�ҟʒ�������Y"PΌ3�(
�/��kJr���o�T�U/�� ��tOW'����ہ�P��>���G�+�%����6m� 4^%!�W��І��QR��u���.�a��	HS�i�q�d�&�6#���7(H�b�ΨA�g����5�>Ol��8���)[��Mu�DbL^�X� *6�ʖ�N%#���L�J�)��ާ��e��6y%��9Wj;G����\�����Gf�&�K86�8�0��k]Ұ1�D�-8I�d�Uۤ�v٪��X@�FY����%cq#4I��`K�a���	⊺��U��aX���hz3m��.7�wA=�$ήVWO�Y�Z�CՍ�U�}#Yw�+��0X���7�ĸ��A"����p�Qՠa��z�(����9�׋��1m+��9L�&��h�ô���2���D�ʴ����Ȕ*%*�8}C���b��h��?NJZ@*���B����C��(����2
@�Az�R4?��4���3���ԫ�2%8!!��Bφ�+XL^.Q]�q����S>�99��
�4�}��fh˚*&$����8P���y˿ܟ�K�$�6�	���=�d �I4m�h���vC$�U-_oP�Mh����ӑ�	5`I1r��z��h�e�N�'��F�'�k���նR'p�%W:����Ư�L��HsA#ֱQcS��m6ݙA4:+�/��pd6}�f	�`(�9-��W���/�A�F�	�7�T�:O򛤒��&�r.�O	mO��|)�Յ��,�@-��?���bK�k�ɟ(,�~���0��aV�CDշ���C"]�zY\�������J���� �(s2j�#�h��'�C;ys��\]��w��c�5-����Y)+����<uˀ�z�9-nɳO��^uF��5��$PS�Q%��0Q�8ܬ ���S�O1X��"Q��Ȕ��ڽ(��T�'j�)�"o��TyA̋���GP��
I�����!M�Wb|��<c��"PkC���$JF���G�{�e�bO���t���"�u�놣���f?{(�_Y\9"@>HT~HX��6x�i�#��Q��N�h�}��
�����vs7t���۲�����5a ��Y�8B�_ل�P)@�c@_��\��,������Tt�8��:�5��H�]2�n�c{u�>��@4���w�	 ����C�U��.R�=��z�H31��*B����샿&��O^����g�;�?�m���Jì�g�9�L&4I��v�3��`d�cf{����a���a�����pZa`tM>��1�_�$���qK�i}��z=~�vbo�5,\��I�v���X��4v]}�^������Gkᬖ�c��kv@߸����G|���҄��\G�����D�JWBls�P�Τ�Vs IX������Y�p���!�+A����`m'r��U7u	?_N�:9JѿYE�&�0�w;�v���u� !��v�Nn��J�l1��.0q�->�^�JԔ�6�f?�i����q�Y��^�2���?;�i�S�bh��e�^�f�'x��� ��_����n��ix-�E �ƋKB�$���C@�MmH>oH��ʖ��R ���`�e�q��'��QXd�Xƭ��C�O'LlZͯ�/��	��O��^pjEpj8��gC"D�����i	�������,�3�c\><l*-��q�!z�d��>�Ym+ڠ��>��eh�۔H!�Ёt�c�R>�E�ڭ�ad��ǧ?�5��)�u���^L/0��@�LX�JK�/� 	^��*=�2�tko-��Y�	�Qf����&��5�Σl��m�ZT��xP'h]�k�ʡ��&C��������v��Z_�k��
|�_ӳ���k�f.����<�%��:��]�(�%��d�4F��H$�w��W6��2�xεn�@��,��B��}hwiM=����8y+��@J0�+�pF��c~Z��ʒ������-�=_�r�B	@L����1X�̬�8�]�<�k"�cg�oƘ)��Wۛ�Ʉ3ǞI��y�Wl� ����'��W}*�h���>�"2�/hM�]8�(�}����l6�&K7\�=ۼ�]K>�X�:�s�)w�QeJm�CTԭ�@�v��P�dّo�>���3��(rf=-{�K4L���Q���U�_��"qdiL�����r�bq����Ŷ����(	]8�5����LpA�/A`R�Zq�ɐ�-�m~b,�L����;}`��oC%���9D��.y��N�tB��х�c�8�a���-������Xs.�C!�k�?!0�]�&��y�P�z7�^AD��rq�V_xi[��r�uٺ�K5b[(��r�@
�w�Y9�����S�,��B��R�c�u4=��k������_�"�u���@����$b�Ac]�C>��\�߅&7��
�vH[^M�tZ��&=����v��#[�[dK��}ٽD�O���z�x)l(����!���N$���غ?y��$�Q���Z��m�Cn
0�N���T�{}�Vr��h�3���7B��aN)"(j�5�?�@��G�a�bǒD�=��~,6�m���^��G��a��w�K�г��ޝf8R�eZ��ҋȷ{"48A}<���V/x�Un#c�=$'Z:�g�5r7���k��-t��#d�:����u^����S�,a�.?��2���vp|�.���ȫ�K5T�1W]2�m�!��:��W_�3��V�U���$�/M�ү9HȔcn����8�ɱ��������u�M�?_�)��)�Iz�v��F{�l���zV�{,�Q&`��wQ���>O��Lt���hclL�O{z��4����3>C�'����ǝ��OB`�d��_��	Q�}Z��y�v�|?ֱ���Q���G�������
��}�PX���v�k[	�b��1ʬ� �'�)��b'��F���t,�	�7C,2���T��`���z�T� _��/�u�滪��T�4x��	�898�T߿$	6K�qA2�lQ�����R���[<���vX��&�CCM�o���F�e��8�Gu&K�]̚��wj��;R�&�Ԥ<]�ܒ?���9�a9-���[���A�Ń�/N}���B��^�6��ზ#͢�ƶ�S����^�0�#MLt��|D72�0,E��/�p1�=����DvF�X+�t<N��{�.h0����W����
�׻��S�s�Á࢞��%Rwq����rd{iJ�%�w��э#�-��MH~4��!����k��e��ÎXX2n�՞xG����,ȗ@��\��9Ii�0Q�4�H��9^�q��*;ihm��eI�iA���E��69Rc�WO�vz)=���.��G��u�m���9�)�'����c�c{6�5ܦ�7	�fR"a�?s`u~���m'z���k�u~2n�f(ґ	#�ej���9Wk�͍��@��'C�P�rh�:R�`x�v��t�� َe���_z4K��ۙ�3�?ƞ����"ÒTn��� �b��!*��ߡ���@�T|���"�*�����N��>o;j�f��;��(�-�]�O�B����LU�C�V/���+q^.H���~~�p/� ;�����~%<�P�P>�ϗ��Zl��>��N�J���Z����V�.т���4�ol�%��xB�����6{Eۭ�&�}�[�����7-c"K��R�ʼ�O���C]2�
'�z���;=5 d(R*@�w֞��٨#;4 C�6O�qj;V)Ja�&~D�)t9�C��s3�������=Cƕ%�a��?3���Cz����X�}O�W���Ki}ޱ��X �WMDe��~vLhr�d�q�r>��lsf�^T�F���4r� ��H�a�6�Y9c�Vj���!(�� F|�EY&r`Ƶ�K��M�B[��M�����t<*���G5�ʈ�-q�KC2l��~[�w���L����Lq�"�[Ժ�\Ć��%]$y�'fɿ,l�Il�~�1k��?���V���'�W����O�2::��]hg@_�(�Aқ������j�4_�h���,��攋��@n'4�Z�݄�Ҷ�t2{�¿�zOE׌���׃�<��l)�{9g�5���X()zv�@�Ɖ���i��,9+P:�ktZ���8��������	�?�M֯۔TU�8�?��[1�bk�NKgyݿJŻY�80��P�\;���(9^(��hNҶ䡔x�����;�6Z�Ȁ�	!#��^q��Xʚ�wԽ�H|g�ۇ~l�V|!��ڸ87w�����A��$�$�d���6��'���&S-T�W3�5��ڟ�
���p�=�\���;O����F&�4=�#�OIt�� ����od�dF�A������Q�N
׷��-F���W�\�I�mr�}s�`1z�b�7�����Ø���w��<b��k��N�qY�z���4Ēf���zH�}�
�3�!` r9'hm4�n]�VR�?��[�̀X��Ϫ�*��|�A�a�L�5{>��{7�^��\5��E(S!����O&n��"�@�
���x�9�쉮�K߁��w���,xY�B����.\��:�fJfԥ��+���d�	����Ƴ���=��g�6>��<jP��GM��/�$!���Ñ��+����Zmq�}�Z�{��'ܬW�x��<�d˝�Bq]��ς⡲ޅ��6���N�'d,�>w7�F$B٧���fV�L5;Z,Ǔ'�v?Y�p��D>���g�a�㖽m�:������/-��"�_p����`
! ��9#�Ϻ:�E�_��*�(?�É���nm��4^�QN�{K�y�gW����m҈ a*[\�eu�.4��|�"�����0Q`֟��ޭn�+��;�ιUDe�:2����s�{�C�rD�bB����"U���G{��y�2�q+��|��-]6X_�̥zY۪�h��9���Δ#k��\ �����x��:�7tT{l�8825����V�o���Շ�f�����a9�A����=Z���.kkh�Df�R]o�,�
��;��l#j���=�g�{=~5s#�'`)/O��.�^U�5��@�4��Ō���(+�N��WKժ��l^�ʣJ����y2�=����wz=	C���nj�$�d6IQy����*�xpJbt��w��
bp��3�1�۱���M6��US W���.p���JL\׃�W*TJ����2�5�]W��䷝������D��Vk��qC��]�:��#f��(s���T4�/�L������X�C�_&�� 5}�m�3��A�������-�?_���w��8�ZdN�d[�[�/$�O#'��2�f�w@�q��M�X �b�ѝ�j��&
��g�M��������R��jE�'Q##�1WC9�$�&�����g)pТ� �0%K�:��|큑"�RVpJ6�B0>p.���;��Q���r�
&��V�e
�����r�G�ee+�%���4�����VH�p�7.��-�hˮ����9�l��v�p>3�$j�tQ[z�y�O���j���f��?�Jl&v����OUw�Ȯ���_���4�������j��ʕ��-����v�`zM;P%�B�K*բ��H`�1����s�a DL%�m���mFG�̔�_�#A���gaN������<f��P��Z2���)0�z�� �Qvnק/�g�`N���clAn��o��?]�s��{���|lt��6��H�������~�;V�@Z݃���/��q�)�W�R\Ѥ�}��|A?�.�5���g��t��/��\d�]��
�����3��y/����"#��Vm�Lgp#z��
=�ŋ%o��S��"�*�A�1�<�n���)��e����"����q�2�KmI��tk��jZ�o$�8�a�yB���;�o�ڮ���*f,����i�P.J;�"�!K�����7b9��I-*Mu'�/�?�6t.�<�L}��c�@Tp���]�wC"�J��Qi��Ol�,���U��ݘ��}�=�2@I��F]^��Z߰*��8	Tq��YugB���tm�Cj q�
�4��7%���x�RD���v`V��V`�ӆ,QqϘ�I&��F��(P,%rI����j�{���Q���1�#MM�ܣ��A��T��3�����bX����(>�_��y��Cժ-�@�'�K1��S���&F5<�^��ĕ�cB���]b�����MQ[W���$���_�W{����cݘ�9'�"^�$�5�Z�~�����T������RM/�	x��[�i4��i��hT��ASC�� k4�u}�D/�r���:��ѓ��yD2���bz|���)]�=t�\(��WU�0����$�_�z�OC�D>h%OhBhsE�q�v�� �2�u��W04�ߣ�ݮD����{�3@L�V �plJ(w+�*i��EW�uۂ+"��%��ՃР�T uJt�F��o��?	���6�H�Z)'~������-����M��ʧ����� ْ�מ�wI=R���z�b�[�[��Q�NK��y�xR��AH[/�ĝ�%ܦ(�㼖��Ȕ��)�<���^�´=ȓ��$��4�&j6��q��A�:�����ʣӲ1�k��Q1
���R>"�kS�*7���L�����X�/����q����f����m��l|��B.���9�IQ��t�R|��puAA	APl�I�(��ݚ�}�Un ��p���f���O�\��"!VX���;b+��r@O��x'Ї���S�Զّ�|��Tc�(vؼk�(�9n�ූ��R ��p)�$T3�� t�W�^s��m�8��C�TӒ;�=3�h�n��Lԕ3�-��E�6�F�� ����R��>M��w|u1:lS��%�����\�sa[�W�i:r�Z���m�Z$� ��A�V4^ ��FߪZ��5(| ����F���Ǜ=�%���g��+�@q����<�&Y_2�:Q��L#�`�� �d�_
՗lw��1�x�?�p�B�В��v��q��ħTcJ⒭D�t���w��Z~�hD�h��3a��jU�c2���`�SMP���a��I�IK�aj���?�ʛ��ꤶeO8M��֫I���o/��z�Ivx�d��=rkma�nY�f
���2�=#�a9�j�3w`>c�e�2��\�3z��
��f$SJ'b�R�r�<R�F>�,ْ~�W5��u�7�:��:���*"����y��]d��Q31Y�n�L��;?8�������8�;7`褸�)����v�stzzDE�ݐs�����V:��|#�=z�$�*�[�������8��dxߔ��݁�G� \��K��T���v���6����`�㔞O���C}��w9����W� 9��"2��v����:���L@������=(�sP������X+�H����]{���=��y�T�"zM	X?� q%q�"�H�ꉙ���Բ� ?F�:�J&WUL��I���s��8�����|� Mo����T���@�V� %��mPeJ]GMe�hQJ�h�QmSw��P�5%v�5��Q�J�<<W#�^V�SG�.��ܮ�w�>U�Q��>�%�'�%
ӧ�/�����憷�\u�?��`���J�=����
�3�'��wƽ_i&��?lĪS�e��n�'0�a��qz��L?��Ig���+�#�����.�R{8rL6�2�7Ǹ�`{6��:?<01�a�� �]���l���̚�C�/'���C�*%,/C����*j����ai����k����Z�Şe���E7<:��G�`=���lΨ�т��$Y��-�h1�~)ڼ@��=�**�F�`�W�X���D5��I���
�柗�����]�)S��*�Ķ��	���*>F5œO�?ٓ9}�	{�( -��ٳj�1�#����������6vDd��oH�se�kɳ`W,���T��X���M
��S�N��_���ZЕ
��p}$��a�X��!&�2������!Rkq�K\�ɲ½sr�I��  8�oȿhr�_8��X�/���F��|6���.K�S�>�k�2��?��<�������MFXo������ e��չl?i)A��^L���_�ф?N���p��|��Ĩ����v.}�D̲�R����R<�Ɯ�I-�p8P���m)�� �܋�c�La�V�r�
=~�ka�����n���6�<���ͷb�k��LH.�n(sI�Uj	}q��8�p�]Lқ�I�����x�2�P�~�&u���R��ç֓
E�-2��r�G�)��<�I�`i'�.��A.�.(������$A�M����*�?��/���k�+��O�nN�њkx��Կ*$�7j���&�r�c�q���Pi��f�eݰ?e������iZz�Tz�E>�tP�4}ݿ	�o[�u/�#h�0���#�K�熯35v	�n�#.�#��HY�}*Pa�ݰ�����_� �N5L�(�w�sy�K�d��6�-<�qS�ξ�(����U�O܎6���>��&;��R�S�6P��X��9M+C�9K�bژe�B� �=2���[��760��n+ۨ~AB�O�����>�&�\ڹOe[:��i/���%#���z&i+�s[R��-�^�Ŗc�5��m$ۆyA^"�`��B��/"O���P��y��c��<Dx#���"�*Z>z�s��c��U�?�1pZF�H�����3��v؇�vN)��{����r����?M���yA/����OG١�Ϫ�(�Yb�H�����}��|w>^Ȑ���U���*�TM�Õ6i��+��X���.ֽ'�;�ʵ�b2��l�H�e�e8���2_�?$���- w�v��&w�[�͜5f��y���T�{TW�=8q+�ŝe���n�M��<�z�Rd�p Yz�(�??� ��u�A	%�w�{��Z�^�+Ґ�ʮ�
�Ը	P��0]�Ñ!䚉yl��< �B�xy'k�\�棑;�J��9��2Ĵ�f Y�(�_P6bR�`r2B��!����Wڮ������*}��:�@EXb*��+-W�b9R����S�
q�	��u��i��@>"\m�咮�y�!�3���
+Y���K�[�=����g�`^��u���QJ{�O��؄����%*8�o m<;�e�3~bvU�U}�o��>����}D�/{������/��iPe��x.�4k�-Kϙ�ۯ��ߤ��Oy�\�/��6{ic}2z$pcK'���%�ޟ#�-�[�,!�RI�2�������0�vkR������	�ɭ�p8!靌fԐ1��x���QF��*�!t�S����� �9�ӏG�E�����q��6�M̘m��Φ�;ރ;�����}����oz&d+�A�#�F?r�W��]f��oP\��}Z�<ǝ��M;�7�J���";��?�������s��-W����Fp@�f�\��O �$=J�Z
X�@|�[Fq�4X�l]P�kلPaY���I�B(�*.��I#����ỲR4:H�{�ډ�};+~�f����r�+~��L����&�m-�������^��DKEֽ[�%��y`���Ɏ�^u]�;�SzT����.�+�$��$L9@��B�=�FزBB��3�R��>�p$�J4���GL���| ��M��Z^pw���0�?���!8�ٶg6IS��&{�ŏ�!�.\K��,:j�X��3N`�]PzZC_#/���~�qшX��c��O�8ᑥ8���\wm��gP�J�y>�">4�PE0�,�&d9���F��j���� &p��S�̀nc!�yxs�����u���R&�R�-\_�Z�Ao9�֏ov��A5��zdJ��ѽ`�5��˚�j.T�i۞@���걫g��w�q��J�$��t�C��E��T���Ɛ�m�P���{�7!Ȇ�aǌ�w��x�U\�΍�Q�k+!��uR����O���(���%0&�JE7��ͦ�I�wx>)�N���s�v)3��kv ��ɗ�_���q�b�s���k��k�FB�2L K�3f�N=�v��]��T�"�!��Qi��c^��ٟ�+�$9Ϳ1���o'���K�j��]f?��oӵ�3�N�O,�����JI����XWB�v:c��zh�V
��H�t�\&ťr$(���̐j�$�v&�=6�?F�%��L��f��d4#B��|���0?;약H{�W��.w/v�_�-N��/�%i�x���N�3�A'�9����cd�o(3�Y��[䨝!d�t{U�<�qԗ+���-p̊��wlV,0"yu� ����7�#����_W<`�{~ҟ�
��@F�x��t���F��	3�
�nٙ��92:}�� �;a��=�Flf�jh�߷� ��ـs�9���AW\-��T��T�.Y㝄���x+8��'�)+qp�,���d
v�Nӕ��rr�̘I�st1��F�?w.��ט�`��\�$�~s����V�G:���#,�ș#� �Ut+oU��x�>�����R�"f��iL�=�+�;I@�|� $)��4	O�x���>��$&�	խ��7�q�鰵�&E��IrF�8VrǰN3 �)��=;����+k"����-��J	C�EHu��#F}hQ����ÇI��t��煣�zݭ֝K��/ΝA�CC�3{u��E�eg�ę������;j|fJ�Q�t�&�F����b�\��m}�8�r�8o�$�`SZ��槳A���ۚ(�o�'�����߳�~0;��Ku�u�J��a�Y�����(%� ���da�7ۋ�{-�se����z3���)�h�V��9�|]��M>&�m��ى'�L��Q����ՆB���sU�V��
������T�j�v6[�e�f_�qS[Q�R�����I�Z�Uy9	C�Q��f���p�Gl�(;.)y�����o��7���!��!���*�d�վ�#��,;%��Y�*�I�c�h��2?�\d�ϱ�T���%�Z������bx�0��$̾�q)��B���@pa��Bi�xQ�]���
��tm|��lLRV>AX)�r��Xa­�!�e�A@{�������V�ሃ ����j�B`-ҳp�	��`N�����WG�^��t��{^�J�I3�72!vڎHE}�濖�S:F��O�Q����]؈�z �)�P��Tzs@�]C6�.�KzC�{�	�m��R �������lѻ���Ezj;�s�bb��{�����5-��W��y�Q�d��b7�n��A��zA�*}���^$�뇾Y��Ü��B/���>9���l 4�o�ƾ�,�{7��:���s����^�.e~�{\	�cq���o�@�0�ߖ�f%)�	��R�s����柇S������`����ĵ�����M�7��o�?@6�-UHmPU|�����H�T�z&�Js�$e-;ԃb��ZG|�lI-�/����PS�r�â��P�3��C� }�<A��h�Q�P3����C�#"��t�y9/�ao@���^��&�ˇ��Ʃ����O�4 i�5df��`�T��y��uZ���T:o%��_����#ִ���s�15��t;�61�$�1V׫�D�2�Ђ��u�����`�f$��y��)
X�H�p�:rnt�����&k�[�k����\��*��E�5�4��ä՘�,�B9�\�䐥=R�=����b����?��B�`Ԟ�Zɀ��g�t{aNa���w��5�5�w Vm��*J��H��N75�ᩄ�	�rj����;I\�����~z�����C2]'
W�ۀ���-�po��T�^�鑂�vo�|S#��8�,�p~��V�,�,g�;K� �k.t%s����O0p��`�d�y��&��ߕ�r��tڵ�����[{��(fu���vޕ�އ#�wi'�Zxᣰ�X����1�,��Z�~\�у��(��c�� ȗ�W�CU���L%�@ƹ�Ž�˃�Ä'I�5��ș�af�5������.6L�Q��X�Ђo`7PR:�{F��K�\�,K6�^��+����kK�nLw�{Y"<TiX���A���[������[��:R�O��]�Q�06t��t,ak|H�W!zi��Xk�1�:�����7Q?�,���J]��g0ج$�'�G�#��V��Y�\ңiP�����sd�߱?n�Hg�|UmAt�r+�,�6���
fV�S�V�ytJ���GA�e��ŝ��5�gd��~2� !�GZY��L�;W�4/�)��7�%�d6��nnF���yAȴ�U)wd����<�����h��H ������G�~�$ޫ��ÕD�-jV�H ls��vi�^�~���ﯚN>:h�E'"���������(�X����t'�O��(�c���@���9��K��hk'�S�T��p�KDI?��c�]�a�p��Z��Ι_8�᧟2����|\�ɋ���i%P�ArN�P ��k����ܴ9O�o�z2
{k!�5g���2��� �F��,��5҅ʊ�v4M $���+�C]��$�Ik���?��у�ȕ$:>��eҋ�e���B����a|/s�0Ͱ����$T:D�J�8Q6a젧�k>\K�|j�:��T[.�
 �i��?!��txB�N3�E�����E��WV*�^
Wخ��h��=��ryS��R�e��6W�	u�X���x��^On��s�p��G��ǋf弖����鯄��Lrq�����u�wg���M�97?�g=�Tƽ����̛u[r�
)�o�G2i�*����ٌ H�+#���ȏ&����\�`���o�r��5���ђzr��3|����gY�g�?������^쟀/��#Ps�6U�S/Ե���u%Y���`�i��oR�G�H���E|a�^"����E�0�(4ͪ��%ڴ�&<�~�CN`�����'E�BY��S`D�R��7�1�^:�{sg�P�[��߬��J	�H!��H�͑��Ad�4�]��;0��1y���NDYc1�49����%`M�W`&O�hv�:5��,V3��\�q؏�����4�]�,S����8���<z��۹��j���?����z)1F�lN���*�p�sTneyRQ��a�+����;�7��UF<�t�N����3�bµ�\m�wTE�6B�[�Z�P\ˌ��q��u��m��~�&A��I{����>���6�e�1&Յ`j2�چҤ����XĴn��U}G�{�B�l��N^�ϒ��B� -kC�L仾��\���4})tR��}J�c�0$��LQ��<�z%KD+�{u�gs6�oJԝ(P�M+'$�,7��� �Ls��r��z��&�U��A�Ά�p���5nX}�����k	����,�D����^�V�^����hU�����G{�)�n����o�H���[�;�O ��
��B�@����v�d�0�gR�l��rص�8�f��d�!W�"a��F�p��=`j6����i&j
'�N�kY��`�.����S���]���O@ �4� ̠Z>(�mv$;�D���O�>h/���ږfy)�ǖ;�<;��-J�%ˑ����fY6��X�H3��r���Z昹�KI�袚�#��%y��h�0Ū:�[�V=���k+.�3҂xzP�ך�UԠ��d��<�$cf{7�\�ф̪�	~����A�o�fU"�v�S�=��̙纶ʁ�>�)���hYB�����Gm� �r�#E�鋵#���w��{�޼t�G3�S���l�qҶYH�/������z,Ү�Zr�4�I��	8�I��^���7��1 <�i��$;|n+|�����Y��$�� ��p��/��'��I���=����K�B��E�~[r|�0�PS����b��7��Κ��/ݥJ�يt��6 �8f�"�F8��g�*��s�F�r���`I�B�������@�4'=X��Y��3��{��l�}/�ŗ7�ё�L�Uבd-B���#��R�ʈ��K/��{S��M[���W�Ō��R��K�N�cB�є3���tl5��=E�A�jN�;�0���Ll��n*,��9�Xדy���m���GKݬf��S�6����w͔����V����>8�ϦI���}D�f�zh��|v���i���	�&�
m�"��?l}�3�)$�f�2.NF��lY�&�m����z�;}H0���j	%�e���ꑀ?��Q����(?gc���֤~1{��$wva�d�?��h|�b(o=�I��3�����" �\Yzl�EQ@ͺ�	!�v@7��V��6����y{#m9�O�{�d����u ���ȁ�ǈ�)Ì�5{��)4�4�(ހ�o"x��}�RxŶ���n)�Y����T�6��;/	`��%b�t[�4�G�l/j��g_�}wdY�x�k���8���?����w���9�eS�+^�-����L�|U�����? #�J-�U�%Zg��o���2�,mwo2�=O��z�>d1�����"v�dI�������j��0���/�Ұ�D�$%1U��[
e��uTf�S�(_���/����rN��-���g��	*��v�mL_ �t���m�\�V�T�5��B�po�݋�@/����!���ž��)/q+�f� ���c^ˑ��j��X*���t�ݠ���'ˣ��g����+�b�,��I6s���$"����G�F�JH�+��#�6|����~��� ~Y�r��P�d�1�J�<�ꡖ �5��n�[0����q�xqcO,H�)�E�"�%���k��L
�!V��ͤW�
����٣{@���w�L,�n=�Xt�����r�q�t��`�Nr���uϝb4C��_.q��S�s��O��_
U2�n�m���z!����Y?Nd��k\�?b���|�ŗ����6L����X�En6x�����&v_�!BM:p�;�0��A*}Adfݩ���'�v�t_��\.�xݱY����A�Z5������TS2m��Hds����&F�x$f�U 7J;>��-+D���2yqP��8�t:�(����^��+ߧ鏗j�Q�'�!�iA'd�*�o�2!�_�Z A�g�v�K.���XY�F��x�VYpm�;#�ƴiI�O�KF!;��c��;
6foW�Sٺd��� }���
1S,�ep$Q`��]<`��o�i�F6�b�|�ID���^:����}&�9
�	����lX���ΰȪ_��} ��Jwȱ�^�2���0��(�+7�t�Ե�IBv|,���J[L�"
�z
X�G��y[X�{�@�`9+I���N�x@�h�	�"�uz(�x,�<=�PΧ���쾭�������s�*����8 Y�$j����r�i*��m-���'��g8��%-�����T��R5�XZ�-?49�Y��[��D����tE��R�t�z;��b%��&�	���+4�,}R�"o }�V?��Z���Ʈ�%�`�sqr��nz��D1���0�	��S��]��:��|�:%b.e���Y��Z�nbS�裞��)����5�pZ���$�2�%��;F��4^�wՍ	�MƔ��ITR�*�� �߳��0��i��W5F#�9�� �����V�_�ٛܶ��A����aD�O�1��iDH}�����§#0t!���ψ~��4\f�r��T{�R�3Hz��4_�F����W��yT0��?q�6I��x���$�g<2>��9r�X-u�/f4��E�;D��
W��yW�άK�������4"�0�_|,f0�iK���ô]+��i;Ia@��*��C��}�����d[�����][t��?h��JKU�N�� �z�9I�#��J|_@�u���׺]�� �v�߹���u�c%�n�|�>�5�7�&E��$@$Ь�.:�ڗ�(ʤ�锋�����n/<W��}VKm+�I��?�y!3Y����)"w�\����&��rP��ai��"�$��:I��`�9�p����W��G�\�f����Ns���O[a�i�w�܃��ȷ�U'��u��n�F�Z��$E������A%&귒%��nbzc��-�~h$o�v#cQ�ք�9�/�=�2ٹ#�i�Fa�b\�es*V�b��crDW	�l�]ݮ��oq�,��^�5:���רK��=��Ң�R��9^=��,({� r��%��^-��n�Ρ"�Ȏ����5�8�q'S�� Υ?N"�n>?T�-�9/Q0A�t�p���}���l���m����H�3A��wvT5D��	�˫o�S��f�{z��z���g j�p �_��R��S��қN�4Ls��j�`rT6���{�z�2
���W�q�?^X=�J��R[�z��1����@���@��$4�N�*���A|�s�YX/�}˾h�3��jˎ�'�1"l����J�
CB}<�*P��}E���>!��K�@ڀ�B�-��1�D��6�r�	�ftԋ������"|�"+��\1*��\*e��{�+��V��T6An���I����5KХsJ7H�V۱p�� �YD�B@��z�s2�x��n�^�4y�x3�͡S��n��z����ؕ��1r���-���oe���?:Us�ti���?;�g�.�r��T����Lw|�G���E�m���9�
�|e<�!�cL�G���I}��%l�	u��ѕ�k+WX�RgMXP��r4�~1�����l/��	�V���h��۞
G����ʼG(
IU�ū��k6j+��pq�6x^xH�V�B�� ���;�簬y�*Ɛ�z�vx��O�|3'���J2l6�Vj/o@���U�V�h�ȕ`.[�`<P�&�{l��$nZE,�ƿ��m�Z��oێ���{�i�-��6FP'{qL�K=���Fo���w!��+#*N�
�R:�������|����5>�wL1�r���-z�7z*.�FA���j�%AIF��e?{ߘ� qP��)+�8J�Ipm]y+mn5 ��K4]�b�U�O��N��`q��(��S"B����ƹW,�?D��|��!a��=뛣ǥ��#����&���&#�|�
<_���f>n7�ѿ��aK69��qF�e��fe���T8��5��f��à�������� ʋetH��k�0R�}�S�����3r�^gls��	U����'КX~�GN�\;�����UB�J�yl<�"�Ɯ)�B�'2�����s]�iO2��&���h��m��M�Eq{NE'�!�5��Xf��ZK>ʽ�)��(�@Kތ���]!�=WѶBb"[��^����;�	�g�Mm�UWq? ��:+TV������p�}}k�Di��@c�I�����&g�G�ox��'��"j~�B�R�h�v��tk,�k�y�(hR�-���!�x��������{�S�9H��N�(�rPC���9~��`�-�ږ��C@���Lm�WM�H��' 3yٻ��rڣ #��K��}�q-pJT�ձ�Q�-�$�B'�$�f<�]�BJ�,�����魟u4@ �\��n����-ce��Vvġ���'ۦr1�b�T% ?���2��+�Ϻ�+;eL��[s��87<��z}�݄ӧ�rbW��"ǎ���;�
1�;�~�ɮz����=�J�Ika���������#b5�<�{6��3��UG���4Z��^i��ȏ��3~QM�)S�����[B��|K�]�}�aD��=�>��
1xIHTՕ��y5�gd���"�,6�UO��}��	�\L��2�����ƜQ�u��H9N8�s5]�ZRtsY[�
�Gh�K�Q
�uKk���vX���7��a�J�#�-�j�	�q�J���5��A2A�R��7]��Et�{�?�Ҭ뵭od�����b��J%�]/�d��<@��!����~�'��c�_Nv����������l֭�$T<��P���k\N��}��?>l�!�ʱ�YU�% &��o\�rL�9��d����"fr����OK�K���n�QNG�ҿ>��\�:>}�i���<��O����RC����lP�*
���;��1��͆����[�yw��:�5E٩���#aO%���&�������=x�O��2j�B���	L�v��T��X�I�{+����o���X`��i����������O,��U<嵊��E+D�X=���*�g�uk��_���צ9i��lԓ�=��.�Z!��������&gb���M������U�����B�NF�"j�UJ�w�x׹���p��B1�͵}�P����\�W��7�THQ��3�3�����D���4��3��T�q�d�y.i��^,�I�n��7e�{��u5]�"��]�D~/�bn1�~��>�3o&���(�0}�=��3���Y�&a�c�Q,�{&f	=3e��k�YO��ԑVQ�'�佶��Y��d_��)��<o�/���9��ϠL#e+ld��͋�ܗ!����d�9�����^�N�������W�.T�1#,Z�T��A4��f7�8��	.M��2�4��5|ã^$m��-[��F#��hT��a\��O>�N��&�;���p�����c�3�5󥒘T��HE�Vs�	t�zw�R�j�=F�Llns|�b�ЌG�#���O{d���{����|�\�>��Ǿ���r	�sxQJ�]5���Laǹ��:�޳����
�3�"�j���M��Iڵ=��.�|5��3/i��Cɟ���~�e��_�%��e��f֚ � �k�>'G&u��z�BtqZB��V��i�A��*[�n�ϱ����<�+�����wD[��:N�z���f@X_F��R\;��|�X X�"˾Fu���6�=�5O}�l�6�z:�a�+�TT�>`h����XQ�V9���{�@co2�_U�R{_]��1��Ly���N��I�<g�1:M؟x�	���l�2 1�$H�3�WE=J{�-�5��|]�<�c�i�$$��lF_�E�?K2Éٶ���Ѭ�zd�ދ:�8���n�r�Vfp�_)�n�yT���Bmh�OT��Ԃ�,�}yb��0�(աx#�z]�>��W�X��R8T�*��ZJ���
H�yKM�Q:Ӊ1�q�H�>DjP6]�+��\+��G��{�"9��qJlE�����[)�o��L� 0Ҝ��U&96oC*@xk����0���'�3��5šLP��U�
���C�"U�X�ȭ���'�Pߒ�T��N�^ZV܂���񁒢"�k��]��;� �|r�jZ�8p�y�%�	�ěT��~���A^Q�K|�Asz�ο +��9����40Yiq.��'��hZj���ܤۿ!d�w��r��oe��-6��J���:S
���{��Q�����d���w����J*�D	�AM���ߜ���&}E
��x3io^t�j"[	Əѻ�r�{�^�汍Y5B&����'���a��0�D��lk�˂a��	�g%��_����R��_��0�Ā�utj�������l��G�!g�W�h�IQ@�o��3��ۯ] �]u�5S�����cs�h�:���������b��zDmN�y[dv�����d�NI�����]jކfC�
�0�#u-I��0W�~~W���&�*�\�<�"YjK�L~�c'bg�-�_7�#6Kba�ة*��4�ZҘ�$O�@	��c�o��6F$1��P�#mq�f�	�~�E뒸0�zI�$� �ӐA˙`�^�G�����;�:�aϹ���N�}�Q؃�n<�ɋ>{:�pqCk�p�ଠ�� �R�:DYc7k���lI�2�ҳ�eKR��>N�Y�,��&�]�*Q�� kUHBR�ݾ��
t�Q�1�>βD 1�z6 �FE(_���;��e���	P��;�Ic!=�L��Ś�k��-�L��+	Ø��{�<�{�YV���|$�|�.�+��[��._
�.+w'~̞���ҡ�-����:.g�[�0�����57����R}��(�J�2�v#p ���9���6��6�mߙ!Y��b��w�o8�e��ʹ�|@}�ĭƇ.v���w�č�}�֝��/ܗw��ŨtkU+ԏ�Z5��]n��N�'TG<CyVc	:�ϱ�D%z�/k��Z���1�x�_�W�px��6�Rݓgi2��7��/䬜_W����1�Іc����"�o�k���C�U/Y��"� ��0Z�_b^X<�)�/B������ }����rnJIE��e=��uS>���E����sW���+����f$ ���s{���Q�#�b��;ֶ���Df�4�& ��_�PR1/�����}�U��"h�e}<� �y`q�#䐼�p�CmA�q��:�lP����s�o���ծil�����J�v�1�0k�o�ryo�Ƹ��ﳁ�|_W�����L����U&��T�TL�λ�nZc��#HQ0ל�O�mIՄ*��`�w�pV�����.�U
Kj�.����TA��|V�ey&J�u�@���$�$����;����8i�swp����	'8��e}��Ptk� I�����X�N�n�/�ϝN{�e`2��H�z}�)��%M G�40G�k��ퟄ�HA���p�U4���*�s;��*��Hk��3W)e�����&�qbm�����/���Y�-,;`���_�wka�/"T0�*
e&]�fu�؈`͟��lIIZf�]w�E����M���0\�Ҏ�${61�|P���9��A�1��fi����")~ڃ�O��w���������j���#f74�K�>�Q�]���ި>�;z��˖NnfZY6H_�ߺ�j��G>�9׾�6T��3a,4������DrѮ����&!=�1��߲t��i��g(�f@ 	Y}�4+�@�a/c�b�g����#;�τੌ�j=U�ډZ<��Hڛ~�p�*�S���p{��S0��<��U���F]~�l�!���!y�8$u�t���O�x>~�n����˰Ui`&�BQ5� ��_'B&pSMt�L�Ѐ�)m��8���0iZ	���:,�o�/������E0q����W�m'�#��jƕ�F(��9	�r�h(x��:i�~�Gc�I�z�H�9�*��ʆ�P�k�i�g�_�d�����u�7N��BZ>�mA�I� �����o�4mQ�I� ���w.xW-����p��U8A3�s��,>6<�v�mM ���*�Z��/NJ�A�3!��,��ɩ������P0�A�\���A:Qah���}K#e�A9C�y�,l`��ຫCm�d�6�W� �)S*#�� ��kv�����k�Z��2[i��!��n]�Վ��FEJ)o�	��{��#/ZP2�˻�[�29�=r��9u-����}��@Pa/P��)1Ba?�	�7���+��k_$�� ˕W_w���ߐʂ`�&yvw�����e�㪬Ϫ���[A�Ap( S�g�(���s2���W����K����-s�/V��o��]7S�g���t���������ﵮ%s�~�	�Þ�����>���h�OlaU��U�j`�t����*�x�������|�IuGD��O^���m6�tA^e�+���7�~�A���{@2���A�V^�ѷ+�%I�kW���4�����������G���3��]ū�j�C�@�S#p���D��N��`���)�p��! �^pi�;� PЇ��<���үܭ��Кy%/E�e�d,���&°���~��x�+�|L[Ֆ�.L3����^T������%-8,kK/���֝kw���܍}%���ƱJ��y_i����^�Q�m|n����;�^`uP��5OL��)�P9,fb��Y�����ZXBk�5Q]��*��(�.�E�w��-�%yDR����!Ao@�T6L&�x��蛒�`�c��V@u_�`0D�E*Bb�*Z0w� ��j8���ܔ"8��Cs�n�U[��������4��QFRak��:#�=�gF�a�]Px�~b�nZ�ޞ�/Ǐ�w�@�2��@F.���vh�4�_��.��K�n�����ƾ��p�:�7�sE")�hƙ\�A���;�zxX%�� 1�.���_q�1s���.8��8+��������!w���lPJ��>�Q�7vjNmG�OkB�O(��w�ּ"1���DP��b8-�>���Y��!�4���j���N�y��n�s�+x��FwdɄ 6}�� Rk?�'�G��Ր
\�#�̩��>�
�xɘ=
U兔�[/̐lH>C�|z�2	�v���	\��ca���d�w����.T�N��G�8�`s>T$��;�R@�n���W�ё����.��>��+�J�z�zs}u�8�B
�f<��]�f�/wD�LZ��E?F5���H���WAz��.��ҹ����4��w@�@�O�T1���M�ϵE��Ӌ�y,�ti�p�j�
o�Se���B�b�!/�5�^�����-X�_Դ�L�4�"�g�s�"jF�e��|�y*�����z*��	�U�2v���2�$���������E�U��R:���̨�voG��H�Z����f�pX��aN�0i�#���'N�S	���4ŊW+:�XC�5���H�uP?UT�*&��A�DAō�y��;�hl� �b���Oo/����FD�916�����Y��]�E��a�>��I^�u������7*�Ch_u/�.�svI�񡕷?(E��Q+�I�z;�$�H�n�VP�S*�+�=���'���@��J���k6ᓕ�58��-�^H���� Y�"�k$���(r�s%ln�h�v眙��������r�1
�m�{�o�)��ד̠<5�5���Hbq@`Һ�m��k���쟦�3B�.�ўCv�f��ot=�O�fY�F@~+n�DS �#+n��X7����wlI+�v���_T���KڑQi��@�1�"�w��d�EX�U���ڃ��ڰ_e�847i����x�3E9��4frΓ�E~]�ɴ�r���-BmS\�҉^�C(�*����J�Y�{�*J��?��Ʃ���&ZG��_����J�y2�7'}��`�+p��TUv
>��h�#*�;-��� ��� hp0�~��O�"���¯G"��E�|~�����ia�����r��7��W��Ějp���g<p�u�0�ŽV �����B�Լ�l�Gs��x�A��jjl�X���%��-�������7��A�i����������r��=�gي��\b��/0��:�:�բ��W5�ʄ�y�	�9��tMJ��`�t'�9^U��r~5��4�|��Bd��#5��'׆G�����ZTa̰��� )�� $f���Iq��2y��V��ٕp$�p�>�L�th�ϬP���u�J�.���@4(�<�U�X��|�mR���
��	��&W����+̹�C������s
^Χ�M~�v�����@ ��%6;��($v�Zr�M�6q2T�7uʓ=z����ߨM��s��.@��dt�1�V�����/
h=��[��\�:�V����3`��߼�2�j'@oW�G��Г�i�N"y�
A*��|���:��~�xv#���g�#���D���b ��
�=��l�p�;£�w�+���wv0��M�p��0P׶A�/�t  H/�[c��($ 
ߴ���:�C�o��ܛ�p�~�LM:v���Ek�����t\�)@�^^���2hw�c��1��7��`}6��	
$w�P"ʿq��e[$��Q[�o�'��b��&���X��N��v-��^��B����P[�K�M���v�z�����Zݙpi�eA��+��r�G8U�����F|�|���>�
_��,W�����%��)U��ÀS��sv�z�K��T�Qj���WJ��Su�ri��Pc�����g��>3��I���˓��QУ;�E��������9kk�������
��7���z�j�樻ϷG�@��c������(�L�f����y�N�5w�_+�����َ���7����)�n�:�1��Xf���K"F�Mq}�R/�s�֭�����Rc��Q�6b-Yb&͍)�A�����]B�a�ŹPK�d1Y*�Yx��-m�]SU�ǐ����"n�v�}M���oW�G�r��I��o'����P塷���Ȕ0��Eq��u����L�2K�@϶���2���g��.�^��X9�r��Ғm�� ��W�<"�����X
orG棒@pHu����$�%��ua����˙�;�k� GnH�/��e���e��7؇xg^�w�j�	**5��A�lX]H��!���THeEO�'�X�8�/�K6��g�E��Ԏ��sG��o�2v��/��$-�%�Ɖ<���I�`n��9�^(���m#�FίE.���\�q}�k�Jy��(#Y�V~�jKQ) 4��3 Â37�S�;�O�F�j;��\��~Z���
��+W������-	s%��F���rp�C-�U~�*�v0JE�eC|�t�5���y[�;b�PCͬ�S�;#���\(����+�]��@�9��e��x�����@�;���◪�袎%v'�������y�V a��ώ����c�P���Q&�U?��g}��	1�M%�>U�P��+|B������ײ(��W)d�7����x�(w1|b{��j�-Ġ{#2�A��c���\x¤�ah���?* �؁���c��<:V�U�e0�Ha��7}O�Hΐ�h��C|����%|�~��l��&#Omx��ر�&+\�s�dtL�9-Kɱ��;�֑���D�&$�{�J�T���!��k �6�1A�XV�1���ֶ�좷�?ܒs������o%���0?�*��*�6��V�.�ď��0����sdS��
����Ӵ��TP��h�L�xYLEX!���ʫv��(<���L?�p��(�͝�6�r��Э�Z)�������X���kH��Q?e�.����@��`<�#���&[�\!q�W�m�n�{�,oМ$��P���꬏#?��E3��pC����2��ID���Q��T=s�o	�a�z�i�G6���pvH��u*o��5Rg�����9��T9���~���W���d�߼Sc�Z؍��Cf+$��O#�� �y_�b�a�ĩ�P_�"R�p+oM�����z�3��Ď���p��'�_��C���=r|	�|��N���0W��g�;��ү����ח�z�iʤI��Pzʵ�6�A4��[�����O4�6���F
:���~@\�I�h���ۮgs���a�8�����rߵ�W-C�����1�)Vî���M��W@��Q�=��A̺�b��� �;�u�L<�.,�Ԟ�ѕHS�����Ž��x�*4���K�Q����5H� ��B�I_�T���>�WG*�T���M��$�5�bN8I܈�M�b�֩��A���+q�^
�F���0(�U�Y5m���� ��4��������ܐ�eA���Mn��� ��l�@��Y��U�,���b�W����=�W���4vOv��\�S�
���+j���D�G���0���<�>��.�\�i�/��c0��Q`(@�v�ng jb�@��v:�Kv�?e�$B#�� ����	"vV�G���IE.BW����A���b֡�XkF7�q��~���������#O�*��
0���?MK�U�%i�o\��𙶏�)��Y�_`��Bǆ:G�2�R^�F
3]o��^#�a��y�2���OW��B��J�#F�`�q҂Α�&`�U�_�����*>Vy^������z{�zГ��0��_�q��R�E�-��k����]���nn��mO�*������5��q��v��`�.����]��_�R׊��b�+f�^��!�ϸH�y��=ȕ��:�Q���5u�G��L�9 )�a6�r�c ��綗��F��7seͥ�*�'P��Ȋg<۔��ۆ� ����IV\�>�4�_Dh6zme[�퇅b63�B
���{��n��|��Ng�u�B&�s�#��(J�l���\͔+|'�-w/vu��
��ͼk�Yl7ŭt�R�^��C�O��۞�=���͑`SV.�q����8�g�\���0.IkW���^\&Rr�֜K��)�!`�?���Ia��*J�c��z�8�u��Z�����j�ﵷ����K��$���4g�_�|�{~h�֔�	�?b@�
�MQ��l�$P�?����O���a0�۪Ez��-�H��Z�������7���t�7�h}�Q?VA#���z2�	i�i�"}��J��b�Ɋ���nঙN]��7� �x�f+�P<���-��f.�fK|O�s
Z��������-[�#�BP��7������ϓ�>�V#T�:5I�w�1���߭Ie44%~��� &>3�9kK��0�����l��o
��)�*ظO��`��L&u��(��2'���R��F��'=����)|	"����!*5P�����eGxoT�C��C7 tYۭ���ÄmpAvS�M������-���E�+Q�))TV���R�uE�y�ۜ'G�v�*������&�=L���}b��)��T�?���K�����#�B�X�`F�O�����x��X�?U�����oĀܖ�����b�Rj˟��0�ۢ����w�
Lt��B3��Ɲ#Tȏ�^6:(�M��2B(,Gl-�)7���b�[��aR�fc����^Y˫�2��-V
D��$	L֔�2W9�Yqx��ٟA.�+'.:� {&��mR�pk}�jM�g��-�r��Ɨ@Q��`P�q9^���ꂏ��#�M�y��B�
��U�p!�\���=/eݽ����%��	^��^g	��ٌ������3c��'���1��X�=Fz�m� ���%���-/�e�������_�7'��۬}w�: �:F��6�9��s��+$wQ�B�d��%xV�)j-Y���ց�m����0n����_�nS�=�RӖ�t�h��nO�~� �T��5ЦA���&?���];"h����?�X�J�&�/Tx#٢�lU���|-��B,ϵ�q��#TC7�
�Br�հ��H����D�\5J<cT�k,�����@@����.J�_�)��ͯ�oj֤Y�ӊ���֢9���wU�T�`��H1��=x�����S�ha͹���NB�#��Lm50 ��/u$�"+@M�()��-8u���jk 5�w�O*��ӓ:Z�nZ�(��|�zs���X�
�
ל���3���� ���
P���[t�Bmkx��s�$�U9��^-dó�H���&|E��i�<P��JW��ޯg7�y��$�jN:�����,���c��\��q��)���F���jZt� �f�VR;ސ]�ӥ뱑D����{��BE��q���#
m~�ذGYiA���]޹��X�gOw'.Ɛ9=���p��;���F���W@V�{�����c�?�/�e���UI
WdP�*�,PF��=`�s�:m��)�ӓHM��͏y������V�ҏ�g!��&�I�����
,��8/��Ȁ��1�[��K?�J
+@8^�7D�gů�K�g�Ƌ=G��%e	n=�ӿ8NE�j$&0��Ҝ?�`��
����?�3˓�E}ߩ��P}�qa+>V���PAu��=P���c<n6�N�gV�_hU!�Y�`1B�K��!G&-����"l;�l�	g�xVTZO���eZ���t0+��S�ܛg �Q���?���Cץ-~�����v�G&90K�V"G�1��]m<�A����*5J[�+�1�&���I��Eׅ�s�"�Lc�Bd�SN��%+q��&�Csg�`)�J��I���O:Y��s%4L�p��x�	o�I���� A����$0E�8ní��Ff;�W�<��),�S>*��5�I|N*MhA���\O�1�1^�}~v�$�����eOh4�$�U��ۆs�3 �$U��������\�z-�{�/����ojޡ��~l��US,��H�/4�̘lkϊ�t�� ��p�K��LT)Z�l\�Gv�(e�^��G�?UJ����U�F��&9��Z�\5�t�����9���6~��2
BU��`�ms�g�?������UZ�����bsk��:����Ư�f��h_.���>~+��
O�-R���OFt�+��aG��k%�Ȁ%�zս��4���ћ!O�3̸s��w�X�<|x�t�s��Rշ"�@=EypG,�&"�n��8ېVʹ��Qh��:_���u�%R���7�v����0`9��Ё�rĂuu����	�ָ�D��'_u:��B�������eE���"�A����rp�*�=��+�����e���0��+�CE�I�h�"��k���s��EL�x����X∐q$��r����]`xi)�$Q���Q�e,=����ڞ�4T��a�e1T���W��L ���\�#QU&�����5�gҜ�v�*�y�F Q�B��|"�k˝������c1�7Z5ey�c�c�A`����	)����T#��4*�`��bG���'.�|:G�r�0D��g3&m�H=ge\~����:�z�9z=������C�s��q��T�(GQ⭉K]��|��1�G�v��%�J�r�0��#B�u�1���`�;��I��C����z��鬢ҳ!w�3Z4�(MӕH�����uN�@�Fˎ�V���Ä��:iO�`����ԛ�.����:.� .)�$4N2V�������1�zYRF������,~���󯌖�d�Qԓ��Y�F�3p�&ݰ90���]
/��_�] �t! l���<`LQ�Au�f,�S4%�i�Z.�\M+'%�2~߱�����j%�4<ô|�h0���|�[w�����C�����a�4�%���Q��#
�	R����G/
é�x����f���=M&�ҁ�������Q�N��c/��|��d;ͤ�I���D8�3�3�?;�xs�x��?D��h�],��؏DZ��* X��fm�KmN@t,$�e�I���H-㶨N��"]]���5.t���e՚�V��0�f<�_�/C�x�{?���,%Cf6��{ �i��i9M�RO�[?���į�0��_���QߗmG�$Y��;uc��6�_|D���2����ŵ$��{��7��Z���4*�p�L�)�(�Il�Qi,�Y[]�SO��w��h��z�֝S�^f 0��U�D��L�[[�<R�S�ﺑQR��]��k�����#��-R���Ӹ��n٢��Yї	�3C�Ёe�/n��p<©�7��J��CjR=�A�[ܑý�k�}S�"�hh�2�.��EQ1�'p\�y���˺��]�7�i"�w$H~+dш����F�|���P}U��s����m贜�,�+q�זn#� �Q�N	��}�N�;���u���^l@P3�bjO�s楕F
ٍ�0��%�,�=� �̽��������w�DY�+o!�Cֳal<���.:J�9M+�|���!�� �BL�����WС���r�Ow��ӦoX*PF @��wȦuw��Y	��)�`N �ɂ����
Wp%,�&���s��Jy�x��ޗ�Q&�Tc<R�{.�6F�*q��vږ�l�?Z�9B�FM~��_M=q���@1��+���ݷx<��x��J?78��5,���@�b�(fx~�r%������^T��a������ӂ� �	-�:N�8���H�� c�b>o�u�ri�j���.k
�qC�V/��;C"��9^,�MIU��4��'��̜f6$�`#+�򻬘�T�����vk�LEJ9��,���]RdH��h;�j@2�g´uXg`�ֈ2�[�r�l<�N=o�9�O�#R��Is6�0>�Y�����؋��^�<�D�y-͟���˦b��[	|-x�n����8u.i�t`���s��0��~5��H�K���I����f�U�D���f�3!'"���s�55�)c��ɹ�MhΐW{>�������[�jh�|oT� �&�d�X����!��^�xsvNj;�')����D���ܢ.�������}X����SU��eA��#":���Hsjɹ��C�~T�\��
��?�)��-�s1�,>y�+Մ�Ѧ�Be%��O�YGCxr�ϭ	^���!q��R��J0~��'�я����m˜8��լ��y.���߶K��o#g�(��utX�j|c\M�������OJ�ℷ�UKN���ڷ�k��NnJ��EXt�S�H��]�z�Ga�M�s����;�|�K�s�Pu4rp�b<���s,�ധlÆ~�[��Nb�ޏ~V9�朿�/�X�9���ђ�O~$ս��t��e4���)x�C�G�a��x����B9���Ձo ^I����`|�G&�?\������YŮ?���"���e�CW������S����@��w��m��6�ї8��� ���v�Z}�R>f��b�%�C0����d�'����+����Ĺ/=�����{�g�Ej��]�ϸ�\d���]R��B�4r;���Id��o��#;O����@dK%�p'�}���,��=Lm��P��{���RS��5�N�l����E���3� ���,��?Up���˱_�f|͚���\�r;��鋪�@瘤lr�jB̢�r�ճ�'s(�f%T�s�a��z=:��3��d,�|�,��N`<L���<H5�eT/6�9�g�Q�IK&��O;O���e�!��9/F��f��s^q^�cX#���p�[�������){կ:���8VIL��LZU�~�4�Ow�	Le2�II�IKet�����u��n�*�q�rl-	Ac�l��A��4�ƙ����z(�����nY�2�'��'��~���,4�4��Ѕ.��vh��<����� ����I�@B�N���t��g�/|"��P��1�3F�xv��#t,j@�� @�+e0���R�J.�"�mw�['�da����%		x?�)'���Ɗ��V<b1T��2L�eϼ�ƣ��*-\f�+:��xz=�|�մ'J�#:qՊ�c
���n���z��Q��l>�0e��������3�;�>~:9s��A���I�ŀ�W�.7�U;�]�P����f�ͶΤQ��!���z�[���̡���(�L^DK�Τ&KoG�88_Kj�@�ϽH��(�]��{�Җ�О5�9AO��[T�k`A���!���mx}��9���R����٩��r�&7�{Xb|Q�e��g�����ӷ�L$��g�����5�6�����N%�C����c+��_�W� �Ծ5p�2����%0׀@o��[r�6
�8�;S3�c�@tm{�4��ia2fQ��`e���٦9z �5 Q��#^�c���U��e�Q���:�'Lq�|�,}!�Oj��PRu�? ��ŕ	�i�Eg�5�2���M�� ���*�M]��F�؈���Q ���NÄ#͢ ��0������%[�[��S��'O&�:&5��fRb�ͳ�~�OE���X�lv�)8���ZJ\T{?����
�1��cK�>&�z���p���`�Z��yk~b�?39��\hM��[�'�ZL٢P�	�g�P�[v�10\�LG������_����s��H�o��F��꼪�?	�\��}X	7�+�PjL�/�EBI�|6����cy���u�"tx	��v�|$:V��C>�\<A*m���4���T�+&��7��lй��a�=oO+�F!.K��5rF@l�"|A`�mmykV�\FP]��!��v,���y�m�p��I�0�;���Rx�w�x�9�
:����Sp�8�6�K��_Yb{�tpC���~�
��}�k�N������H}3��$������l��u�
���2݇�*B(#{�?֎��[�'�ި���A`�u�\LI�PDb���w�/g����l�V��c������`���Aڤ���u�(�)�Bt��t���8#�9��$8
:�D�\�^'}q���L�)~�j^�F�(�c��!�a�)�QQEТ��*h][!��tɁ(�Z����4�sɠ-Ok,���ٶ�Qg����JaH���/��/�������Мuq"$=3^����DT�\�c@���	#Q��y]a���e��RD���	{��Q�CR2!��pR�q}�x���z�C'~���o�Ԉطq"�j����;a0�v�v?2��&4����e"�(?������>��d.��ܱ������Y#�� ��0�q/�,�JP�`��=��W�_��5��5������lH�g�z����L�o�Z�K�Gc�=�R�p��n��["�5�UQd$�=0�h$}y�'Z�1�0c	PFac�����>,�\�?\,v�ƳR�ДV�l�9i�bҴ]�b�k%y�la����e�'��#3`��^�Y���'����mˈ�a����T�	#��v��t8��˅eOd_��e�G��6��b���sq�%�Gy�wyI��|M�����̔rk��}�6-~�#?C�N�5���zu�Y�H5<�g��Ih���2�3�O@̵�	��v���s�ɇ��'������Kw���j�ݻ35��7�0�lF�!��lzb��wz��]��3���]�}������ A�"����������(eI^�#V[�w�7�Ը�R_�P������%,�b��8b�N`��Z��]h)��Y���*?L�䆱�!TN��"�:����z��_XA��埻��H%[�̮�&Rt���x`(+�l��y5�Gt��m��&xR���f2^#�p�KL����w�RT0�"��xA4�u��q�T.ާ#���S�Sv�������4vH}4�DTI �-�F&Gm�~�V	�I>��cDɚ<���M��M
�h�V-���Z[m�bl*�p�mN��"��Y��>�>�Z(_�X�D����FK�GP�/3��V�J���|�^�V.��O�y�݂�M
op-�o�J�H����e��0�g�mU����Ms�f�w��T0w�۟28���f��yf�!9�<��"��h���[ت�{�g��>�� �e[��Xܯ�Ӻ�Dޔ4�F��*�;��(w_q�>__����}J�Jr�}"ᑍtN�v^S]6�F�|vʿ%)|��`���Le���֬S0D)�kPxQ�y�}9�quYRX�ytu^G��<^���mÃp�?���V{��kd��| �Wz���h��ѱ�3���ǩ3���\�o)_��q�AD"n�U��XrB+O�=��׏�[��R��Q����s�!�K�I*H�j�'،G���� pO��I��W����h�F	�x���s1����0&�����İ����x�ox&�|�eМ��7�C�̮���ke�|��i�sv8:�;$XTb�����������R�����1��2+��t:AlF���v��+,���h&�A#�#2��A��ͫ��GpӦ��&A!��!���n���/DIo�v
62��2s�5�w")e�׫��MK�n���.���A�ZgV�*���PL�����k�a���cO�8_�Nk���'���`u���HVm�\B��jxA�y���z�'ğ�k�F�d��%��%��8I�,+"��ޫt����J|G,�{z�Ec���������0����jT��&:ܭ�
�>V���D����u��A�e,D��R�g��[ԯ3�Ǵ�p���0Ff���XV
;�w����ye#M0��1��,�������2/������
V���젗&�������+R����+��� ���a�h�%������4P'�O�� Q�"Pn��=�vs��JUBc .}
"m �����2K�B�:��w�#`�>6O�?ǉ7�K�����rB~`�-^N\Y�6n���6�a��R!�$��������I�:�h���ΏE�/q��P}���WB���U�j��d���c���&�n$"���4zI/��oaXIǷ��5{}�O��"��f�;֧S>���_w�fUO��[�*h��������TT�%���:uK�������i��6���t��� &�$R��-��i�$����,Y����k555Y��/�"6a�0 �ĝ�ǽ���ђᒩ�ھ�g�#��DgK�Yo�NRk��C�d���B�g���{d�؊������
��v�~R4����b�a�M��?�P�U_�L�b�SbX%j��	��e_{{��`BMV\�w��T~� Lc+>P*r;Gx�XG�˓�E����Q�=��]�.����j����K����2�hG�Ip]��mke���~R�\�����d�Mf�eEtD�E�̟Ա�N���[�<�S�D�:��3E��j��Ċ�8j�P��I�H��\04Rp�Ю]�!�N��s;GIgЏ��#b(�Y�j��<��TJ�2A����YX���FD
�B�g&�{���,�F�c&�4)m��a��_�� P���DE� ��\�Bkf�_ ���"��>�������ѩ���11�]�� "9N����Sr�{M�]���M�k�W�'�F8t��(8�oy�o�x��Au}c־�f_�ɴ��8�h�K� 2���;���p�=v�U�/�m��jj�$욈�d�SP�u[�D	
�RkK�7���i/�\v�$mqdaʻͤ�~�Y�T�]ɡ9�y$��y�b�1Q��x���թ7�U侪��2T�J0�����P�r������=�Ԟ���֟P��`�s^��֘GOQH���0?g<���<���th>N<G�C�;�C�����5�n��K�o��1D�\�֣���i�:Vj����
]���\���J������:8F �M!W(���R����x���e�b�'t�1&~u.�D7�Nb���� �k@�P%/� ��KXd��O4-��:ݴ���F/�k�ه?�Z-y�,����H8{�.�3��zqB�E��i��CCf�JHY��}�?m� ���.�����j������!ռ4���Edf�"}�k^Q�B޵lL&c��eT���*/6p�ߦ��}q�A��O|�)��[9��\��t��X_�X+\��,N��Pwue�|��)�glc�rQ���	���t��A�]���0G[�=]r#���=�vWp��C@�D�`f��H��H�]^���r��g��`�i�C�z�u1����Cg[��]/��MO6E@!�m5o.egg8F8�Om�9���yѬ߈I���k\ &n�(5�������n�U�Ҟ6c(��I��Y�}$\�4Dwu%�EH���T�_H�feMV��6���v�_�I#=�kb]�$W#^��k V <��%4�x�Y8��'���\	�x?;�h#���O��>n6��1�7^�\��k�L>�[���f�$�����m��d`��	�q�&���k�^A׫���CT����x��Ib��Ǒun�7F��#Oz���"�^7�N�h���Kٱ�S���HX/������8X���^��fby9�Ĝ�VJ2?h`g�kBl*X�4�����v�P�Xu3��W��1�������x��FzfY��s5c;~9'��#dsqS��J����� ~������쇊ys����囵�7���z��<m�YY���}1z����|�Y�!�Mر)E�I��/8���8P�0���aW�n�jŁk��/���-IƽFsϟ� �r�M���Yüq�i0�O�b����E��(�L�9Rl�X��e:��&��]�D��Q���G�K('�� �q�~�q������{S�%����x.���5�'Oڰ���\�XY���Y�2�C?�2�.hf���z�WD���E�pV���'t=Æg�8�חq�}��S�@9i�"�ـ��."@������0����>R����T�ȋ��h�Q�O�Z����u K����0�����Q�A�6\�����y��ޗ*��1�[�6����-][J4a��J�zas� �t4�΄[RO�~��Tlu��p`=CX��};(fԜ�a���l=��Ӡ���yU���?��{A�5�k���	v'ɛ�'�"7�j���zs�?�t����J�x.pKg�
%0�:t�w���^����n���C�쵝�K��񑺢�4��2P㞡����c���s�wZ��1��̗�@����+�1n��%���S��>��ɱݼ�i����c�Gڒ�k,0c9w��f0�Z_͍�$#B�����<1�Fi�8�^%�&]�7l*:���*M`����`4\p䛩����tn�B!
+�BwR�*@�1ȝ˽[��xBT������7�Än�/���q�AZ7�<�F��gU���!,W��H�lMYʦW��v�Q��6�;ڲ��&%��t]a�TBݍ&����B�����1�R��9��W��p�X>nuz��) 3�@�ns�ǽɂX�~�={��a��zB�����Fr&E[���*.�2���x��[v ����i���9���jk��ap�"� h��?��sd���_�pJٍ�rװQ�T�x�/�fne�-�Wa�bzL���,���=���J��Y���1o��â�8��S��	�޺cH��u�cD�z�j�w Rz}�'�얨�/0_v�owҐ����f��K�J=�l��K��)Y�.�$C����օ����Q=T �q.x���+6�Jh�֨>dC��z����`�e�Hi���������sB�x�%���cs*�"�	@Ⱥt9E\*��hfUsP��)�ट��
�\;�f�W��;�wP0��԰}��8y�aH�[-����E���W4��7����.q�����[�n!��MbE�f�8�0}:�R�h���;�}7Z�UW�ߋ�?jΗ:t�~��_di��HΔ���?�5ȷ���C$�8��ѩ-�so�{�e~{�#�W��7c|`�YWJ!, ���������A�Ga:�ݜl��Y2N���'� �v��eZD�0�I��̦�e�4�יF߱��X�Lu�E��u�c�C8mE3���9&]��m�Y��J���A��ˇ(`>�4��'������f�Cg�G��г������/���FG62G��BU��K\C%A��E��ȱdt�D��I��]
�$p���_m��x�?;��nӟ�)�w䅌��"Br�B��+�+����� m�I-4ɶ��#�~� \P�e�'\��k����;ª��*����<�[AVw@Q�_3Ó��8�y�r��d8ۄ��O�Q���U�o��X1����Z����#B���:/�$TVĤ��\hs�A��M���PP`�v/�:��y�� �<f;)_u	�9נI���Ǣ�H5�˼���L��c~��<1XÁG��k��N{o���<��e�ԝ�i^a8Hh.��O����P�OfZD��&!�5v�����C����7۷�b�_�G�����V��WRX�hgT
�RM�~����\��u;жr4>h2�(��U��總g$�3\��'v���z�3EN�3��.{�ߪ����I#m�(��)�iR+��g�E�������pd@#B4Re�,�'H]!BPJ䛣�U��S\�6��`W��ߩ�Y.w?�����@�?�YR�0���VM�L��>�����KSn�%����_.��I�Lu띐'9P�_�m�勺lO�5�/�f�
;����o.� ǁ����9'|���^^E��6������:Y�-�����ř�Е����/�`�����$��N@�5�t����o?lY�y	Ճ6'i�6{��DdɋV�X���<�K��q���a�(w-UTt�t�����K"`����1��q���>ߝ���B��&��Q��u'0_�S;�w���aJy��	�{��2�c r]��,��F�����t*l�,��*�X�۠&5s�P�Ĝ �|��gɘf���g�E��yn�-����\[w�2#���b���+��}��)��UL~�MMR�����|��,D��_"�Ⱥ�t�x	�ܵ��<�u��5饬 �'���N�j㟯Cw
�G:��sD�s�,� 	�4��Q�:� 2k�@/ӝ,*�[׫�����#'�Q.����j�
�5}���X�a8��-��M<e[�Mj�ԅ��0R�"ǐ��]s�a��h���"��r��WKO�����0�T�l-?^M��s�-t��xr�i!�Ĭ.b�'6��z�4T�8�����+���pp�M���}�'�3�n��	U:*��3�;�!
i�-�A���&�E�D�u��k�����0�$Q�)��j�ۖ���I��x�!X	)h�����ѩ���ꓴ9R8
�8�k����X���LU���O��xP��rt�}}ٻ/cZxzl�MgG�*�7\;yw$+�:Ӷn���7��|��L��	�r�VLK��?��m҈���>w������� n�����d������Z{�BC�,���J8;���i� ���I���_�?Ԡ�~{��Bmήv:;���`��/ '��\.%�O!�͵`�ڠ��E��;���=d�[ȫnCYRƹ[oР��u�ܪ6?N��6_�2���F���O+��H�ϊ�ba@B��J'! �ͿG�$�!ϥo�fi8��`��� ����.�̟�[T�k�?JNd��N]���a�.��b�X��V�JH��lǠ� 4�_[,J�N��}�j� �ۺh �u
(oK�!��p79ԡ��:6�^~��T+] V"w�x��ǖ�m����7^k�O����y���N�|@t}�`�u����J��r ��Q�[*{�����!.�������O9�Ӽ�̈�NM>4�i�A.�o'�w_^����~}���1��.�A�t<T�0%���9��j�+����-�&�$�9��uN��4.,u��u|��^;d�u_��s��>-<Ͻ�!��5�o+Ӎhj�v(��h���� W�����RH�Dڽ"׀$K��mI'-B~g[#W���#��q;�QͯY�s��uo&�D,�>.���hG�ƈ؂�eF�$H��q�� ��m�_py�$��'�6��<>��E >֠�4/�y��P��
[��"u�W(���{�K²Gr��q4�7��@6	�UB������>L,6X��H��E�ou�O��}��虹$�_}�Xxq�,8:��vL�#3��� zj2�VHy�v��h��*z���l���ޤ�L�=��y�JLEAb�l�j�&5/#'i!� ��a�yM�K�Ab�}�C��ur ���9	��aB��1��e������/L ��}�vy�s�J�$0��,�� 
�Tp�c>�����P�5r��`��8}�ؙ��q�yO%>�#~�]�2����lĶ\|I�ec���ؙo�Dz�Q*"��k��'��i�g�<�N�򤼸-��w	8�&:)MU��J��{�k!n������x�dZ˴[$t|�%�d���m6N=ٽ�@�^P2����yh��r���k�{8����;g�!^����8/\�h@�.=5� ̔z>M��ce�q`����|o�k�8���ݚ�ǝ��3t&_b���g*7�'7�&+���F�+�Հ��{�1���)���Q>�8)�ڔ���P"T�m�*S��r�${;m:����^�hv�Ut�qa��2�e+��!3�̐�4l�����c�zDf~)W�	C�Z�M�G;e	Ԓ�o��ĵ��O��/©��ȥ+D"�sb����{O���L8FӁ,��֙���i�f"Ko o+��z�}1f��U$��i�x��L���r���k ��o5�!��gB{�(�D)��+�34W2�NC_]��{k˒�cH��,	K�0P	'�Uc(=��V�<�`S$�1}ȵ��?�az#��G�̓�{2�:���Z^��+VQ�W�Ұ��H��X�=�W�Y�9?�ǵ��:��␒�/t�l����`���U�B�W�[Un�L���ރsF�m[]��}k+��w#�^a%���Kо�����󛡙1���9w�0A�-��(����ҝ�tC~��P�V%����f����{����Dm�}��b����ǛҰ��1ZQ�wL�h̊S�qЌ���I�i���Ŏ+͊]�Ƣ`��w@]��3�Mk����P�yA��\�U�Pt!7����EO6c��^��]e1�i��0�Z����@vb4d��_,_hȨ�%lh�:R��#~���V(�ܐ�J�l�~9��T�Q)�~쫏͒�)x�^�x�Z0��/��0�x��\��ԃZ-Wc%i��m_مz����л!]�X���jkֱ�ң`Su��s�u*Tnr��i���[�X�\W���i�@��<�����zxK���\�4ڕh�.�!:�t&@����R�,G�����+u�]2S���R*�2m]<�3;��()����G�#��:}��RJ<@.Qs����~L/��z��tY򠍫0j7���(y��� �}���� n��(�q<4�M#�(��{�� ��nJ�R��z��a(T�˺�7�����Kpe��h�
:Js$�۾�_��L_[ ujP?�8��K�]���0�~+2DY1�.�I��ɳ��+�)*��>�L8O�l��w�fct��5�)�^�c��mڴv3O�����W�!�B��i�S[j$����N�1%���l~�?k$�Tˏq6ؿ{rQ�����
�k�q|���۟QY		�@H]qg����;]��*ą�9������]s���+��̾�9�`����Y��L�CC��YP�ge�a"1����;sU��>�>[>#FJ[�� N�٘I����.4"j�}��6�ɡ���N�� ]Vl٣�Y�!�JF(����G��i��l��r�D"¨Og
~okT���^�5�ȸ���^�৳j8H�h.�:Vm����jz�g�̭E�e�7Cj�˖���7�n�N�$�h� ���!I����m���������Sz�4���joq|�"Fd�闵�`H�;�o���ɟFU�|&U�����?kE�ot���Ȏ��qg���M���M�KTk�>�/�V�]D-oި�ZEc�~ŃK9<o
�ZI�,��8r��Zq$���L_�����}��bRQ��邚�ߒ�����f;�]���<�LDn�	wsP��"[�7��A{��4�����.�#R���%��rȏ&}�!�~Aw��W>��ry�l��X�W`�������|g�����iuq���)�۪���ڟ����B��N4>�[%����z�|��k�ū�^�-_Ş�����]<H��m���ۡ09�:z\��-l?´���sDe�I����q.wG�Y	2�L;����JY^��zW�2�#ml`���(�؁FX9Ϭb�_�H#���4��xf�B;����>����)o�ύ�뉯cKOB���K@��&��Ή��=��(:��aHS+���vH��<ڗ"�?q�f��^Pl���}e��?0V5X���4�C�&����tE�,]����:o�5��Y�'$:��.�If��
�du'�^!�o�%h�nQ�����f�ӹ!&���+��p	��G�+�(�v���x!ȿt0���*��@mxf��5`K�9�Ɛ���J�Cҵ�TGN�G?��0�P�`�w������T��ܓʪ��,��͑���L;��:���j{��!���~��Vh�v�x��ts�%�6J��A�1:׌%�t�k�`��!��g:���DM&k��֏��F������ h�Vg��W�U ���i��\��>�H#�A9��_�#�%g�`�@2�jQ�,F$�kgU���'��|�����Ui��R�_��9Y�^��t���܏�$6��:�;{t[�w4Y&�=�^�?&T �dQmд�еr۟�s����~ �&C�W3�x+YԲj��2+DD��s\�ry2��#�6�r��X;�I���D��H���o�s�p���2��DUB��$\��`�Bʺm�\��0eAbƼ�܅����{iӟ���b��nWDT+
�-���}�>f��+$c��6Zg�Oj�>} 	»�F긚|4,���1�n�77�k�z�3���A���|�H'���P"'�:a
�N�-�����g���R+���vabf-,�۰.��&�x��~��AG9�B����5�e���Ll��ڙ�͈�:e�^
C���R"�(�:_�k�=R�'��k<��(�f���}\�mn���Mg�*Κ،'���:Qܒ�ݏ����0���63���2�Fʶ����u)ZP��@Q�6b���Y�>��>�թk�m����6�0ﭴȫo�u}Ewﵾ���͈�C��ѫh�⺛��9l��cf���z�����x���.^+X>�	?Ũ�<��a�J��Ija����K3���}��o�N��_5U��{������Yc+�6afd���g��t/����Q��HD�����G7�	Q�@��:�ё�ӌ����*Q�(�B[���*��}Py,����V�xb̴�&��RY:R/�p:������tJ��H:A��P���0���	�q������F)݊��ֲ��T6���ewJ�l[@��H,��ڊY�ٔ$�U��N���U�~���DpP�q�Z�:ܫ�}�qx�n��o��O\� ަ?��?���{i�A��`�ǖQѻ���J�Z	�a�J8'����v��FS�H� Vi��V�{��g8 EWn�d�݌��Щ�{���Zt5���r�p;J�(*��K>��w�@����W�sҷ��:��p�vxlzT*utO�f�*�W���>��7�V	k_i݁FN��2�u���gy��TS���M��w��'�-uƞr��F۰�<%���1�o�g�較}݃��J\�מ�����.>� t�C�s_�*`�J����:�S2[�&�X�	:\R�^�$���Q5g O��"BENs`��&����uZ��-;_�"Jc�C(�>��~��U��i����]9��1�2�Cϯ׽��˱40R�f��B���?����l��n��i��`�Z�bqR��d���1R6`=�(��ڿ9���E�/�{���������3(�x���
���?��^֊�f�Q+lp��b������B�{���O�]�_������4|�|��A\�@̢���x1�e�.�UIp"�_�0���_�>��Q�
����gQ:b�K��0��n�8!�!��!2�r����R����g^Tjװ��c���L��o�ZC������|J#�Ɠ"��j�V)n�Tӊ,m(%/��6;�:`ه� �G#�+�C�?1�P�9c�%��'Y�e����v��Bl�J��'�mAI�M��c�?���os:��$� �nq%1�yG�G�粌�o��a�l x��L.�c��*���#�3�����R����6���Ы/1���F�N
���T�͊�c1�@G���@��1P�p�;5�c����nF>b˴8#���\�Дf  k4!�8����bH��4lI| �:�c�S[m��R��7(����D|5&����5�+���>Y�.��X��ʡ�*�]�Pwti�s��k��� ؀�{����LmcM�d���:����{��(gK����k�{G�0�X4�,
W�#��M��va�s�ȹ�ć�R��Z.@A2o
]W���1>�����B�������c�Ik`МqOc<���_f=T2����::�U��;0LvB ��
�/ͷ�e��O
����{ � ��~zJ 6�y�U�� ���g�LB�]c~Q�R٣vߺ�.���i\Řɛ��1��t.�6��e�ȭ8nZ �.���RlD�+�x<D�/x�d�)zd:ͦV��tM������{q�s?[u@Lَ�뇬��bL�WVq�m�״���q���m�E���C���..7S�nwxI�岻���+Y8�DӀXJ�&{p���ؑR�7�ܜ��+9L��u��ie��5��,���`�r�M>����K���6ǧ�b���}�\;�������ԏ���ȧ���ΰ����E���i+O��o\&��M#r�r BSF-�����=5Il;�n,^t��I�f�V#1�;��-Ǔ�I	ưp+�	���qW�'��/!��e�?Q��FC(�������4�E��Et:`��~�k��]6xv�cx��|��x4P�i<�5h�¸�V5�usIVo�e�/뭸M��Y�I�#z����4v����귪ц���x�`����;�]�p����,>��h6�ٵ1nt~�AV� �hTzs���
D���6{�[t��#gg�6�SO��&ȽB��rm�U���x�(n}�^������'=�=S��1%��������j`'૚t�����;#��j@��eh���z_�|)&���1C��z�2��}��'P}������T��hz���t����j%���h��li&�)^�x}+&���j�Sg����9�Ep2}P�S�����p���Rjp󭅀4b
�-#H'm��_�����t�t^�А^��tLlST=���f
���!/�>q�q<�3��iq�x�:"~C�(Q���#S ��p�us�x�vU��葳*���5����P߇���
E�Ez�3�B.Kt"�$O1>����h;5Blc���rW��d�7��;�A�k±2�ݱ��RQ�aZe�{�OZ�X]�bɞ�AO�q�O�Э3�b69]eH��ĸ+fW�d����D���y�"���9я2n�?���]9����(��W�uX���WF�`��"V}��^���h��3�n���t�fh~��UE�*g�f��.�&PZ�p�GD�oӡbʴ!�[����i��J�(�b0M�&�~��ղ����͌�ּ��{'
SWg���Ũ!L(�~��X����E= R���S%+�JXɦ\��+|P������َ�Ʉ_dDs`���˖��@,��@2ݏ�v�$�|0�ePHC�4�M�?X[g&� Gɡ�B���e��a}np�c?5���j�o(x�`��e{�o�ЖRC�+`XM�A��le�0w��5�jA!�^��̵�j_��J"J�%<?���2m�k���g�W�F�_�f�]�Y��
)V�R���7��M��e�>���d��NA9�A����Dr9�#,,�2��L�\�T�*��=��kw�����6f �^�o�>���b��ʊ�W�,�����$�ڔRe@��]��s��7��DDcg�^ 	53��]i�$����?1�W�+�mx�9���2ݏ�;�k�5��*�y!�"����_���hgo~�zY��]� �;]�z�iV��aC���Y8s�0����[�F�p�|������q�J� �N9f���[���zk0��\�V�SF��L~e�s/��&����*`o���Ϸ�O�k����Ih�G<�*�S��J�x�ՠ<C�ܣ;�_M��J����?u�G�S��=AS�e�١+��hW�Z�:^.�����1*���"J����4�sB���_�X�1N��|3w�}#jP�r�sR)�Qс�]�ky*�H9��?fZU�Yo�j��Z\0ۏC9���:�N�(����Y�Z�#���Pz������ ��6�JF���bѱ�RVɮ��'l: ;�3�� S����/��IQ]������MWOp>Y"aSO!�����Y��4�q�2's��kf*i�5�]��xX��4�l�۶6�P\�8ӋNil/�� �d��$�K�Q!�D:�{�����L1g�}��K�u�߂ϑң�Q�`>m	�P�WwB�X�����vN�O �MƇ\�"�(X���A�h��lw�ȼլ,�^u���4y��q/��)>p����1kϡ̪ģ�v���C�bw}6����+�� N�.��_R��٬�.��'�$q+����i��t�S�^��I��d*�VG��4s�!��u6TxB�k��&mr=�F.��O�L��lT�[zÌ��g`e��r�� 'h{����"R�� ��l��呔V?�]��	��M��O��ui&1��~ ��S�i�ƺ���X�#�RaZ�p�ۮ����yp��P���1����=)g�X������Џ�8l۱f�5�>{`A���i02]@cS�thvgj8���bVl�5ǁ�����$��V����e�\n��f�CZ�Ldus���@�S�B5�h���Zܠ�ӣ��à�h薦Lq���� 8vUhRVL��hT�^�_���ȞU�N�7o�>��}�2Ё���&��1���덀���l��vH	��DW>5W�Y^�0OM�׌e.�~$n���W#WG���0� M��{y��+s��H&��D���mV��4lG�]��or�N�Q�x�Z+��f�I����XV�ǻ�?�y�����f�EEe])Dfڀ䒗�wQ+�Nu{f­��=|��B����t)��pB3Rg1�����iZA�r�[)Y��J�{�ų7[�)�g0 �>M��>�9q�7�4�1X��Ƙ��M�襌�ݼ�!s���Ѯ�(�,�5�b^e������ܓ��>�F������bѩzG�J���f[�^O�����aAQ��1��P�Ɉ`#q��. �;��{�A�O!�r�1��;�ށ�kq�l;�d�Yr�cyl~�J��=°�����f��O֣E�Z@�*k}�l�Z���ᓯA�o�7�g"��[:�!��{�a!-���a���
���~�+�{+I6�L?����!{JѶ,s�Q��ݸu^V���/�k*/��#�!vڝ��O�|���9�R�z�`��غ�R�#$�խ�Z\���댚+؋��'��� �r���u���aK6�"��ђ�J��ti�P�׶P�JQ�b�t�ބ�-S*aH�W�''�Ѓh
w���~���YKf������������U���_��-z��y��[����hbN��E�br����] ��bޘ���F��U �!q�eE�=����O�m+j$s�_�ݽ�`�nڪL9J[���{x~��o���@�U�6�>h�zTԽ��-;Wˉ��G����0�:���C�Q4J|\��Wt�W��^�7U����f[y<J4�ܼ7eEV b]�^�(���ݓc��*������7h��+�X�% :Bv��� �<xwP��t%i�y�y�����˟�E)
ׄ9��'D}rb~'�t�u}���@]`��9��zgF��0&�ٓ݉���?�W_B��6����F{���6Eo��9�����ӑ`= Ї�X�^a��~�5l�.ڨ=L�M�x��zNP�MB9�g�׆/�Fn�y�B��"���}<].�Ǵ�l�S��,�z�V��^	��W}F� [�Íџ�j^�Y�T=m��[P ��&��hS�|պE�t�x�}iH�c͡��x*��h��d%���+�
��A������$��E�@��e�P��Ri�i��zC��P��Q
��-����7xŀ}U {y,�K��|W0��惸a-��@i�ZT΀?~�da��������a>~��8� �6���ފ�|���k-/��[�,f�ռ'(�h�j9?�ʷs¯D�g) ry�+5^��=Wɶ}��p̀���?ԯ�Rc�l���B�W/$y���>�V�3�
�T�H�ȧ��%�5�wn�Mƺ|�+����r�?�xF����r�/�&��΅\RxF�_�0��6`6t�	՝�5A�m�UF����+�YR J/ܠ=�����Z��{k;�54]K>�v�Ǆ�(^v���x�|�����$�
gSh3A��\v��vCA�MW�MJR�©$9�Ӱg�� ��'o
� y��?)�]��(F�`�]��(:�b��s��6��D��3���M� .����bXS��`�eŅ�RJ�B����ˢ��E�%l��wS�!��qm�0���\�Ep������'�>N��Y[�۞��F���d���ʓ H�4'�r������w ������^��Ie˔|�ۦ�'YA��A�ZP�T\�� Е��{�W�`{J9�HSC��
q�R��i�e����9z�?�mp��R�cu��C+86�û/�����β������Eb�#6�B���_Q�
��K���a�n����?H��dz�Jkn��ƐvXs.sq���L�&8������/�*a�惏
�K*˵�\o���q�� hn��_ '�=�;Q/i����6�jw��t!�������w8�	�����D�?���2�n<�w�� �����<�|,*������j�����������Z��0����+�#n��%��mMNK���_T��k��F��+�}}�����F�*vú�1�L�(8TOU�����
�T6���悉�.��F����<4Y��x�ϝ��� im2%�A���;P��a3b�kłϱ�2>�Vl�����_E9��%�����K���G<E�؄��5T�M�"l*��Y�0�ù=����L�Q����I/�pw��es3UY�-|�L�"���8x-J��Q� �N���QC�,_���qS�kJ�T���M�S�����B2H����'{��6z-.�U]�	Ra����"���5�&��Gћu�)��Z"��1�JTkR����w��rKH�lP|��L�ŷ��4>SX���z��2��`ۖo3����!�+?�?v��=�W~�Q|��2��s�1�iP��N�������s�v_� c�`�M��hم�P��*�E���UYq�V�M�y b���-\>�>��3��1��a(r�m��q�}!�v)Q6���D(s�\�!���[��T���m�*�g&��B�Љl�i���lz-7����h��^������۫v�\WW��!e��a�Bs��0��c�Sf?����N�Р��0M�=����\������)�SZ��$T�+�tM�{�t#���7�4��f1b�&_�z�� \�zMFf���f�#b������{��86�������-C��1������R���P�`�}&���k�4^���� |�����ƹ�j��,�c�쥎��8鬞��M��`}w�?��_ڞ1��ҥG�����,{e���%�z��9�¶P�Ȯ����GB��%'�R��ܪ���Y���{��W��G����uɊ)8o���#m�?��kB�'��m�0�>zW���k
*g�!��Y�Y��<�tw+�� �������b�T&7��_��:7���'ˉ�8�Q�	��b�~�mY��v�ܲm�̒gD�ĺ���`��)��U���P�U��R� v@��n�!�C� ���z9J�*�<�`C�FH �|-�}�s&^w9( ��5P��$�a��ː%Hp*��$L�ܔ�T�X'\o*�OM��0h	������-�+��~Kw�iu����.��
4�<J)3��>A+C�B���w�T�U��r?n5�?S)���]ž,5^�E����#���#mD��%21��dǓǏq옰��B��s\�.ǆ|����Z���`)�����5���_Ry¶
»��Թ�>�p�I�]dƳGG����0��4�i�C�X�<������h&��Rşx��5ؠ(�ͩ}���v�{�I�����6�"���d�Σ�1P�\����%�'uAp5���%"�1fz����F~��=.?;�ip��h%���D��A����F�6�]��Hĸ��2���>?'�N3t�m���>�|t.��<���k��,���q�C�����%�GZ�Q�4<�S�D}�@\x��#�
��P���/����A!0X�ˣ��q>N�� [O��S�`��g|�
B��d�?��}7��i�Uj�y��>x�kE�vI�s�+R�����Z����BNn)Q�M=���'?�C¤���s� �=� ��v A(m�L�+FnhT��Ny�a����p�������uwQ�*/ݨ��	udM��~�� �@��k ���טJ-��d�I�&Z�H��҂�{#)��R1��u���M~�|$���Uc1�=�5"�zK(��G�t�x�:Q��}/I� o��_��ѐ︂6H[���~:�@
>�,������JPiZhnRd�&qN��5�S�-Dda�����%�{s~�m?YB�O�Z_��;�Gm,umԮ�;`ݤqd.=G��P�%��}-��av��N�ck_�ˣ�c1�=ˣ�/C��-7�Urn�Qg��^�O{[�@����j�c�\���I�v��j=i�&��]a� �SC���=���#M*N2�^��=#>�|���;��a����KJ��{�L�S��H�g���L��W�]{c��N��k��^y�������Hp�8�~P�k��3�̄����>Fg([��[VN�T�`�tS�#����*�9#�x[T�LF~�Y>�%���V+H6�����=7��N�i�͑,"�s�f,ٍǨ�����Z���?i�h�A��]c�?N�r>�j�{l��R����'�Q��D61��ݝ������٨6���Ll�7�G�����;ȥ羟�1ZtF_��Z�����5*�Bc��ɦ�AeS�r>J�,�g�Ҕ����7��.+��
#bU90�N�7e����F1�b��PmYSҳLN�I.-�D�.`յ�L
*��9��1�&�Ƥ>�	</�wS;�>�I7ށ��b�0N5w�
�r�r�"K��S=D������s���=��@�4$�$Y�O��NY�-�AO}�1w#l*-��&�c���S�&
ก����&�Y��Lm��3m�8d�$~�ϐ�%X��_p�@s�{�Gu�M�SS�p �'lN�Zg�1�����?�ӿ@���ELh��޹y*��{��������Ѽ�?AH�Ƨ��Ў���WF9����[|�c��d�2 �[4tŴq��,0����G��Z�t��%y���Yr$�}I�*�Vy����I�ƺ���/�/9l(�:�s���"I���Ut�#���lW?,����?�e��x��U�(d�@���U:CM���DZ�*�?B�q2@�9���$�?7V��>S��g���,%Ձ��2����^�^z�~�]�a!��S�i��_/����c�G�H�{�\$F���X0�%��zgz|� |0I��� �!xk�/�Cvߺj�����4)`ꎦ�t ���]�~�t�oD��B��W݋�Na�����pNp�U�)9u���[է���(�z�9&�}��V��6u���"=��,�8^�&�A��9ȏ/���;k��ܛ:a�����=�����#Ԃg��Y�`
���]����I�35� N�S�(T�p�"�F�	�����fM���q�IU��>��]Dٯ/�b�Ti-�1����2�Rn
I���d�%�#�Su�{w�V ���Aaȍ�U`�z]�]��<�-cu3��ޠ�_8�xg�<��B�d��.��os��}�ֿ{����ә9(��dj��hC|�l���3I�P���0�RI�z����T�O�^-� �ܱQɛjvE���9�.f��!zv��R���Vfь(�����I���Ә�ϻ.���'�C�*���6����)Oݖ���%��EZ��A܌t��&UN��3K������UK"�FH�~=�s��b���D��F�T��M䖀�q�J���hہ� �޶����䣱��E���X��||yߚL]1�#!���	3Пb<�I��j�Ƚ��"y!���SK(�)��6���┛�%��I\�� ��_z�/��קev������Zj�Э��O��%��f96BnݜmN>]4ㆌBǧ=���̓b"_����3;�04&=h�WЫ{sSߏZ��=�5F���d�r pZ���#&S����"�;A��ύ��SE�N�5�kKI�ۂ�@��n�ɞ�a����b������\�-MKاϔܢb^@j��Ɯ1��#�!Rc7��ڗ�ЪM ��1Sѩ�&J�Al��0���I5�s��	�,>Ҁ�@DI
 6}��b�>��6~8� ��L�n#Lp��jVzXj��r�J>a�A��id"o�8tߧ$�ԞP
�@��'����������e���~LR�(ioy�+}��:*"���|�~X ���)�p��GHG��"��$Y�[e!�Fb����m";"��x��6��53��m�w�)�4�s+���n��,':ҡ���p�߰-nF(��ck)䐎��h���м�[[�ʮdи9@��,�AF5DU�Jq��)*'ܡW� '�^*RZ��5���FH/V2+a)m�
S5��.��᮱�φ)�=!���)���\���N�`��9xߐ��*�ECX�c�wN|<b?�	D0P��B����Yfk��@&�\��o16�]���P��%��{4�;xm,w-U
��M��[ҁM�{��Djۛ��Y}��v���i9����wn��{�����B��t߬K+�B$,ψ;����/�k@�Sd�[��/~rE^�Y�a�zx-,�������vn��$8p��GH������\�#߃a�+�&����(���,i���W��B��9��cLC��Wt�`i��L����S��\=>�/ p�.�uYzz;�krg
�L��?��Q\c�@���&#Sku�EtZ+��K#?�I�7�`�h�g��wl������U �_�%o�yh���RS7�D����&l�̶Xޕ�q��s�)��|5x��K?$��9�0Rܡ�Y���`�n&���ƯFÞjo;f����}4������B{�87K�XgQQ7�� V.��ZN �59Pө���|[�а�>�Y�;�0٪K�}���� hٴ��h�2��ř�w�%M�2tĽ3}������+�k|�,1Ic��k#D��}�Z���O���m����c=�\hn~�J�):=��m�ۧ����>6d���n��Ɩ�U���񟜥��#-�������<4\"��5����:wپ�F	8�6��M8��$����m(�;ߔ(��-QU*��i���Ґ�R�%�{i/c,¯��Y�^@�������7��.���͛PRk�>��a@Q��/I
WWZZrC��
CF��������a��Ei�d+�!�cC�[��A�D���d;C�b�[w>oH��j�lx��QyS,�667*��VJ��D��S)x=�#�*�6��%K�k�i��c��uܢ�u(�.���_!�q~�t�Ơn=�YO�q�X%o�����-�~�����6�����a?Ǘ�3C=�i��W�
�nD�~������P�)|Rju^!;��>c���h1WB���~��j\��������;[	m�B��!݊��
�yi�R^ �)�kd�I�V�9��ubag��]�0���p���$�=��m�)��*FI��}�VukTl��ASqY���[���ք���;�/!��ޫ�9���;��I?���HYxo��C!�6�`ک_���1C���Ù��Nƴb1�Wm�k�ԭz�M*s�J�Q����RS�5$X'j�}�+��d`�����~�I�#���Z�m�G�;�(>�Bט29|��3�l�	'�DΉ}E��t:v���Μ���P3�ڷU5���a�ܖ��_��s);��|�C���ۍ�v��k��Υ�0|^w�����-����F�t�'`~��Xd�[��9�����#�2�x�p� 
c���'�U��uR��S]-&(6���B�F�tXH�iLFE����J8�"y���8A�n��2��=�}��6����{��>��Х��2^���@= y��X���!�����.�v��@w�&t�ygǻ�Ý��Mq&M0����g��A���ywU����E��*#-<m�O��*.��W_w�Fu�}���zJr!���^�ZD�"l7�� h���D���jC@!���|�=���k&������HC�������BEl�����J0��@Tv����h!�d�`s=���ř�s��*,��{��\laVk"���������ln�b9�9����Y2(�[��af�����nv�'��3�@:�2W̗ш���c�̿���p�gֆY�!>�UK�6�{yF���ZC�S�B�1�[�.���D�Z�8֣�$N��W-�2S�i�������D$�ŃPuUL;K����}�6�w�<�:�N^�5��)�2w*�m�/y}���`U)��U�.�@�k�\D�|"���
�{G-��]��q�حwG�k�ٽ�>R�c��ݓ�oK�C	����.Iu�r�8�t�? 1ǼT�Go�AM��;�i�ȫ�a�2��V
�$��j�"�2�/[f��y�}���sTe#^o�s�2��5��@DrB�r�	�3J�`�N�_i�{%�x:��POn�
 ��ݹ��m��j�>��&�J��0���n��ǲ���uS�x���6f�P�?́ &�X������YP
�i�U��`�\H@lE4�.���3�ĕ:�,���Ng��u�X���+XN��2>3�:5rꁡ/i��K�ª4��dP�a�p(��Si<��3<Y�溋~��g�,~#V{y�a�Q��0PF&�������B��/��Xk�d�y��O�1E:{!ڏ�G͗���s<p$��������v��VG��Y;�$�e8g	������ػ��c�fG뾪�!�鸣>E�G�p���_�VB��8˂�5Du��}a�.�*i+�v|��z�H��&Upx<,���/��^�4�34}��bbW�h����Z"i���H^�$U���s ��S��ţo�I9��3$��!\�\��߆}��i�i[D���'b&k�I�UI����ky�*�:��2#3��m�E������
fb�k��`8�C5���k�h���� l[��(%f��7] �m�c#��"�3	{�����݋`k��6R��rԷ�k0J���&}V�&8ʸ��!/�@���ɿ ���8q�����>�U�P�%�ǵ*X6Ki7��[ϓ�� ��]mA�q�kcx�*��b}���x����(#����	�z U\�S���%�^L����C����A kp�'K�fq1kZ+lK�T�<CBY�]�D�k��\U�Z[
����M-nF�r��9�Jk���W[���Cq�c�SI�"x�P�|�j�f�ZDOn|
Wr�0��P����fŠRΈ^�.�W&�G�C{�L���0�IT��)�r�Zc�J�+OU{>l�ƃ�0_0�j�[n�!���]-$��\ 3�Z�H�mH���J?���Rq�B�o�S�h���ۈ,q_�y4�3sw���:���mn�H��C#���hz�[�g�FL��S4���ҷ�öd,�c-.�ԇ�O�&"ƎH��$���הߘ�(��=O��4�V�a�p,wx����!�6��� (�n�aj�8l�h����Mn�$i��o��m�6�l�
s�S�}.>Aq����kxpq�����%�5�f4�[&B��-ʝ>.���^�R�j�m���Ӵb��)���/ ++���O,��Z��Z��������a�Q��ѽӓ��s������N�"է?�`�mhWv8/�=� %Q������	�0ڈ��x���Jo���ȼ�}��r�3��gMR��FT����޴3hR����l�(��&�~�%�)Yk9.B�P%_�&$W�9��Ǒ�s�;��˱�[�I��63)�/�m�p�F�Q�z��@W��NZ(J"�]F^�.�����ka�QV�ƺv0}6�Ll�a�LR��D�o��c������<%�6��?��^:�J' �b2H����ٍ��;V���KU?A�"�_�-Z�P�$훀l���7���jys̚W�H���/ 6AT��,�^�s@Q��g��d!9ծ9X*�f��&Uo�Ek�b�-�j����8��2
���S�4����r?�ն뚂8C��3ǘC�_�jThYEc��b��$r�x�&{��u��Ӳ����]�Hڋ�{��|�4� ]�2�S�	i��^�a���M�#�ث�4T
t��-�%���.G��І����S|�gx#g^��Q6�=]�;1[.��-Ψ�CBQbb�Z<�&�+,v�ȶ��������ދz����Y��Ì6φ�E����b|Һ�<X�
� ?�^S;yZ��ΰP��)����4��f~�)�`,qc(9~4��p�"س�cۢ�����ҽ��.O�-cN��TTy��h��k@ ���!�J��`ėR��#	+C%��2>dV��,Y���5�$k[Du�:0����@����R��*�ӣ�@q]׀þ+��̧yI�z�krA5֬Th өzC���l	wA1�Xl;q�
�meL^�Rx�| ד&�0��;AL/xk���?������$���U��Ν����ySCf�kJ�L�W�"��<>�f��	��9so�A�zꦎ��>@���桑NT��eE���}�X�G%E�co�JdKW�c�T�7D�1���jC�qg1���BHXn��~lgԗ�~��%���QPm�<����c����r��߻IH�U����wis��r��bTv�'�$��K����a�qw� ��)�U�(��>f#8�h������k���t�#�P�Xi�8��|����ѩ�½���!=^q��\�������B�];��)��[��.�?3��ڔ�1��J5O	��a^�z�LTE�RG|����^�!�yӕ~�ln����O�����(ʤu�*�YW=|Q��6�ɇ8�8�T6h��>�T*n�d�D�摙����MUi�;a���oC+��4�`:��Z�L�Cc Z�=���"c(d�D�k0�y��fF8g��u�N�l74x�ɳ��;аw`�RFM��}��:�!Y�,�_5@�w%:��?J� �۹�N�'���"��E2���"IGY2�]�Β+$¥.%�����6~��CE��XKVZ$�:&\���Wo���X)h�o���w�s�����0�y��4�ר.
��t�"N�kᚨ�@���]�
)~�[<�
T����L	9��z�B7o�I?��"���f����ř��g��M[���{zv+u 7�NC�}TNDO8@.�pZ�����
�/�$�������b �{�-�z���v��`	Co����g`�k���'�~iv1*ΐ�F6���'uIO��ZMoAk�����~ɻ�
������P���m?��V�	d^A���މL��W>�
SAX�B_B�Ӯ�9�6싵��,��I+��:�
�Am��a�͈�7H��կ=��Q���ء������/B�ʥv1nzR�h�>5�J� �UU�S~�vKr���i�&_%��<������y�qAp&��呖k��Jy��jf�^ꟁSd����z�����1/iR9t_\��A��Sv7����z��ڃ�Z�Ʃ�( �M�f�T�/� ��ْ���X7;�SYL9|t�����s<>��^`�P~u��%q�������̪����s�,�� �	��f��6:��ٱy�����A��\�kE���[8�D�[P:�t�I"9\���^�Fax� ������QG�Ô�T$��=���w����$M����x�P�d�N�:\��M>Lȸt���Z�	;(�~�w�V%r�=p4P��c匈���w�x�r{D�������V�VF������*�Ǒ���=W�*I�k��6��36J�3U�)�@�^�ֹə�!i<(0�	κ�G�:��Bl�pn�*jOI ����F��C�i�
���>:��E��2�w��^�e#�?��/޵*\Q3f�5�'h��ʕ^4pO݈��mԾ��I��������l�G4�l��-��>�TT�7����1,�9��7������
��ߑl��S�Q��
`d��N4����/��_K����щ~9�~R�+�9��S��{U=��[Yp·����K ^V�~y֫�P��:1Z�,M+�t�����'m��$n$G%�u����� r@��jP�R���H�Ӟ�������t���q�^d邅��W��T��8+�hb�Ւe�7م�s��j�9�ܑ3�� ��a�aX�]�q��:�4�j��-�.�a�sz΋��p��gM��+�;���1]/�3>�>VX=`}���zQ�;^��h��XO�^�W�(��7N��hS��C�,�8@�]DM�K��K�ʁ͸,;u}5��}W�MD�޹�5��G:�ͮ
��a��)}U�#nO3��!2�R*��Ϯ�wħ��MoM����s�2�M��k�af��7i�%�#'�k�K��,ܛXF]�,s�r�_��%Zp��
�΁�r;��u�=>ܣ�N �k�Y�����[�	�1�ť�.�	��qߣ=���(}�,82劙u~���M���Q}�����[�?+%&s��6��u:W���נ(�R8+�V1o�SH:yd�{+��kk�;�|�0^�D�4	{[�W"�GG�㳛9��
��,ׁ�FH���]�k�
��"����:�(<LQ�� W���EH/S�w�x=a�UY+�ϺN�1��*�@�ʣ�bh �$��↵ �-�39D�1>�Ԑ C�y�ڐ�Q�z*e���E�Qe�|mv+c[��P�����G��yvSB^,�T�����Wl2��3��Y�;��w��W���h<:!���?�ex����'�`\���m�o��z�o��{�@�n�D�q��{�͓��N���^(�~�֠�_����[���T�\�U��!��9�$V��ґ�,6W[}4� g*ݳ	�L{���
��k6T��P��hez�<s�G��-���%ӴI��"�'��TƫWEXA�4��0Xtb�����.�j�Hr(6��F�ю��Hi��G5�3�}zmQ����ܐk��w�)�k�>�l���&^k��9��A�,{)&�c	6���pET�*1���A�!L]�5,,�5�4f�86�%ɗ�{����t�&��2��Sf��
���E�;����%kab@�lK]�)�w��1/��m�[����Ge�>3��<��^�a�L�ܨ~���	�֞����1���9\*6P�t!T:�I�o��$����4*������(�	mI�M��Ȣ����u��,j�M��z/��8`߃w�p�Co.�YW�����g_��|'�B��L���+���'�ܿF�&�f/�2�`�RD	:��xl+���K��&+��o��RYb��Q�tjf�,�Yga�8K��8ysԐ�m߄r�s&`����"qr;e�t,
�4=��]T��0�j���Z%�ӢB����Vi���X�ݼ#��<v�u�34󦎽�����[�AL�Еtǂ�̽�:O�J-@T�p�hN�8���B����743�Дϸ=��1�A���/N j��g�����J����֓�'�-t:)�'���oe���+{j4�s��ݰe�(�0e!i*�b�ϘЌ�?�vX��,#h*c���6/>���	����B��.�G1aϨ �Zm�y�s,"���>
Ԗ�:	sN;Х"���5Z'�K�\K��� 1�ί�t!��EAԺ6K���z��
�"͞�F��Y+ �N��������،*�T���Hل��V�|�0�Zz��1�ٯ �z�bgm����21���b1�"I�5��s%)��Mډ�����m_�*l�Ƒ�\��/���4��d����E����L��hx�(L�~�>��wڦ�|B���)b�(q�	@C���욓����N�t�K~C��g7Q���Z��.��8�oO	[�r8���afC�����R��� :��1K_�L�
2��/�	�qʼ R�`B�i4��ezm�	��3 ���pU4Äl�m;�8;	E�K%�w/0�2�������ד��2�Ϸo���PU�4�1��1��V�wg�&��O8Q6���.{���&���HK��9jx�g����GX���{��^��Ê�z���zyEw�c���~��]�������Uaɑc��X��g�4����iZ���=��FNc&���`o�J;�J�ص!zz��Mܷ�^UK[2�~^��La��c��ݾb����@�C8l!{h�4��H����a�#��| �:Z�Jd�
g@���9dS+`B�WrLM��|���6o��|�y˚2�z�����Š��qa�=��o�U�� �R����w�ǋ|��|�ځ�˿Z�1���v�����{>�:���-ϒ1e�Ȑ��<Ĵ^	�IҪ廯�C:_�1�&C>*H����)�+ޟ`���7g��*ґee�6�-V�D<�[��w�[��:(�(ʖ�mu�H���DCm��L�Kv78HdDO��k��՞��bZzd��Hy�7�䍾F��KO
�Q<��g<e�b�T�zw�mхW.��ո�ݗ���q0	#c�r\q8��pd�{6���["})|W\q^J7N�9b�:�^�@cͳ�ܾ�#�d�~�7�
?������ywNV�]9�E`su��X7����늞�z��°��z�&��b�t@�s��-�������4����YW�词́@��$rdl�_����7v���n�$!늄mC:xt%��w-�; �nd1K�ѥ�����x�{\n)���y�5�d�y~%M��9��Y`�'O����rH��~�o�2μ�6Cir*����z����a�
.Z�,O���l�ϼզ�M��cبE\Ē�t��.��)a�i!f�:�?��l�ȵ�,�i�PM�v��d1*�б���+��ĿwX]=��6���+�<d~Pİ��1h+�ܫE7��~�'}y�^�������ఫ�1BZ� ��M�H��װ�6L��vywH�?��(��(��O�UQ6�*kez�pu�����Ҷ�#�ԎsJ�ۗ�~�Z���D(�^��A�Vtϓ�(�f'8����� �����V�|��҃��L�7���D�q�Y�{T8��'����t��J:�[���cpqפ��� �pq�9�NH{�@�G��q��a��Ą�~k{������(9u{�,L��wy4d�OS��~%��p�����j<#��9�G$�-�,��L��v�=���3�S�s\��nN�<B4�@J'z�r��|��bd�_�7�y����c��.N�5{��ߣf�/��ud��ül�� A'���
�A-�ō�.:�S�ue;�8d_�b�ӈ�$ �;=�GT{��N�bA���:�� F�6��<��S��m�w��cK�W�ͣ'0���,�,P��\$㚺_)����y�ϣ��؛2�*o6�HP�&����v�נ#�7`C�������eU'4/��p�
���l�2�<.��+]�����t:�V+.�11N԰ �ŝ<_t�x��w�7>]�ᛖ7^���h���.�]��
�j\��$N�ƅ�	H�����o۪Rw��H�ҵ�\�=.G�K ����VW�	��ظR���ρ,uS��LM��T�r�������{��<���u�?���ۤ��<��E�U��|��_�ٵ��6қH�:�8�L�\�����/_Ç�Ɖ�%��p�6���ɦs�%:��d�艎�g��t��):6���)�X���g!�K��T_)r\u?�Y{5r韌� ��""�on�����[�e��峕2s	� �
��G��K���TҒ�/����@�?�;�<���$ƛ��3ܚZ�ӧ~c)'s�~�3� Ƴ��A=�Pj^�6H�~��dq�-��J-��MVM;M��Hp�����9���
Q�.�8�Z�*��O9wk9�(�4D=�IS���[=��r��-
�LQ��T�-�BD7��Qw���$9! ��s�k-7��י�e���T�|ed(g�L�-��CK�n��*LFe����4���ߍ�DNiMl)�(��
o���0U��o��|pA���$�C@I7��G����v��������E������I)�����`�:F��
�w%�~�iEm����t���A�K�"�2Tt(e	1o_0���W��	�� �x5dʊ�;Hz[W,9
������������A����i2���>�����W�D1���-ىVmP`�ȭ�?f���qC�<���Tբ=�Cl�.hۇ���������"�2V7��	�$����q�5;l5Zm�m�J�s����5���U���Jr�"��K���O��%-�Dۣ/լ�'~Y-������{"c�S�|;/��+�A^:��]��E�l�����>>���Ql��bd�'���I�έ1�'��N�[$]�p�_��A�	���DA�n�Q<�I�P�ãP�TF��K�?:�ry`R
�G} i#�$���1���)߷m>�nw)[S��
�5�-9iL�#>�E�H�l���R,c߫�+>�.�,�`G���� �̒�a�:ႝsf��q�CP�n���Dt	�r�`���`���O���Z�r�� �j��2x �*Qc�۩y��f�?ݺ��!i��29�~̏9?D����g?�E���m)��iō<�9ݭ�4�%��*�!��cy�`ħ�6�,J�0�h�5C,I �ä�i����<,*��QǇ?X0ǃ��9�Ė]�4kə���]s�v�T���������e�կ]3�oߘ�}��v����&;.�ǭ�] ����,$�h�J��|L7�}�+$�#b{g��b�˧����� EX����6�������b�Z�����������hZ��d���(�1��9�G�s��J*F�������������m�(Ȩ$3,�z1�o:�"����V�,?��fʷv��+t�JY��'���;�>r_Ĵ��j�:�h4YPY]��Ef|m0��M�s�g�@���aѴA�����p��z�G�`�+e�����esʚ3}9�8+t8&��/$Wy��IKgIN^h�c�׆
�p���?Ve���@ю='I���B#���4���'��ڮzK��05��O֏�����zK_�6w�R=�_r0����K�E�x���S�fI���J6!vW�v�pU1FW�9��u�)����h�H����Ű҄V��e��kN#k�5�IUoRZ)�����L+\Y�#wJ|�.y�����qM�:�݈OӦu��vB�{� �ww|oiƾ���R:��vSG�v�nB*/��x�̒�0e�bG�"o�l�����T��� qD^��a���{�p���[O�>�C�����.�Kq�%��A���+B��ѠR6;F�=纠�%{nS*��0yv&��;�̀����X�83���(�h0r��+%<�����B���ŏ?����,�[�=$N_�\���;C�c���� ��"�;{�@���m��������4�l��,A�;m=<���� 4�_�L�V���E�]=pm���E�j�忩9t. f˳��J�&x�Q  jB���{�����t�����L�6wo�8;�Y��(�;W�5���L&Ҍ��KP��<�i�N�D��w�8����nUΝ�Cp���;�m�V�e.��
J <�?=u�=��2�m�zg7F�B��#�ںb��{:fv��[]��m����Ż���.|/m���z���@OL͎�56[�6�`R�3I7P�b�J��ɻ�I�
^v�"k��pZ5|�\������L.k���#OD�,*G� ���
��e�~�y��Di��f
�@n�z+Ɩz�/�H���8;����U�)S���$=��Q���([��lH��N�J-X�!�'�Ta�E�E;�G߀��p��ܙ��_�-O;;E����8��$�٪愥���.'/���5sHq��}���h�I�Ȱ���<�.���	�
|bO0�m�
CJCo��ە�T�=��աv�49OB��(���q�=['�o�<��b�Zt�t�^K3��Ż� ��w-2��Msqٝ���h$�N��=��=����%��Wk��+���0�si�Ch0* U��6��:N�c�9I=� q��N�*e�|�,�F�z��y?�$ae=����xvRyv��QPE��~~����M*�q�+�]��5�a���,q�����5�OCXdRɫ\;�E%ِ�ɗ���xS�\V?�8ņD�h��0[F�/�le��&Cbʉ�����OS�I��%]��pC��L?C0�Dd��.��~:)��7� ��19��B�x0�nJ}9,�������+�*��W��ࢮ��Ac�p�l��:`yzht�`�غ��@�b��S'�y4ϲ!+>�P��Q��;�8u�5䅣䯬C~�Q�p��f2���f����K��XP|�Al:�m��'视�/�8͖<�}O�-�wM~)���Ф��� ������jp˙�"WQ޽E��1N���`Lzƻu�bL�d���bV+~SJ�:�Q|���HH1�0�_��E��;+{��O�`;߰�],��G*SR��cL�gD�����m��3�k��6��e���Q�^Z�?LC���i�aH��3Q̩���Jr�	���`��?��b��r�"]��A�k�g��X�L������)��z�H���'b�!^ZL���6���<F�AP�����6�3?��������w�.zd,j"9��L��)!p����I���-.�j�[�΂_��U-�5��}��y��������4�sl��a�(��1��Nd������l��s�̅����&���S�#���ފ�>Ңz���H�-����}�""�{94��L.Il��7�`��
	7��u��Z����Lؒ�d�n`��2���:���v��&�]���i��r����}#D;�9���?�v�Ig�+�of��w�]��jE�o���tg���١0�SX� S@��N�3����0��k(^�,�Kz��ye)q���&��M_uќ_}��VVL�MyrL?pH�_kItƸ�m�N/�6���4�j�eZ�	ih�jz��no��ߢ�$��Vܓִ� p���'����7x�DBA����߈M���M6(�b��Mp����ftR��h�d���T���*W�8��}N�2X�:T��4�&���Ԛ=)& �d#b�Y��@�z���
�`H��x�^\p� �0Ձ���yၙ����xĹ2~�/���8�����9e?Bڛ�R�����]̀��5�@�p[���'6�&�BR��V���V���;���D�jM�Ԉ��¡{�]#W�S�D8���!4��吂`Pe�Q����lG�Ы�ʭ��s�;���R�@���|�ă�N����)���T3�8�ƼX��y��W��r�R�Rj17B�qx�t��F��71������_��G�>��w�3�e��y^Z���"Q���N5*B
��k#��G�傤v[�vf�p�7i��y���g٥|�%wu��+ ߯�.�s�~��I�+!獊D�JU�Ԛ��I:Jl� N��$�>fK��\�|��pEgF���'$�9t��qpt�ԯ�<��y�3Ը\�#Ig�P��h��o�j8>�[7F�#�+>]3Il�ο�kҒ��Gy�����K�P���=d6!���+`-uDXoC�l�;���)��9�2o�8� �����%*F��RN ��|����w�ۃ/�&�u�RŐ�5t��T&#�>/us9?�^���ؾ%�-7���L�,�����[��/��g��(�1�|�$�:���?Z�� �c�		��i3�ݹ	�p���XNQB��o���%i��b�����4�Gi��x���6ϔ����,��Լ5%���j�,�2��;��4?f<r�2��×1{7�&����=_�����EXx4��Fޗp��L�`GLmX��ɻ�W��!���f��Wp����m�@�	齝�2ȿ�-z�dnA%��-A�h�+)>�Ze�F(���GgQ� ��Fk<|5�]nc��ڸ��+�0�vJ
�r;fb�$m���R�k�}:|�8QY�>��9�C]�uj ��y����E��N�-�3~�|ź��Od	2(��W�V�AI��G.d�68�S"��~�2�*�?�
�DR��tOl@NW̧	@�w�ϬB�z���g�����G��l �Z��b��j��AP/��e�9��eO����0A(2��%���@�X�+İ=*�!�A8�<y����rm�����*(�4m��m����������bt�v\Ss0ݵ���-��"��!�?j��g�k&���q#��B��EG�'�	7��v�5��ӯ5���25�g.8�2������?y��2���[WS;Ǟω��1����U�n����M�����RJ/7U^��WF�Q-�`Jv�s��D���;���U���5)�F���,&���SXj Lr*2�"�0�6S��oN��?�,�g3!�~SP�x7j���'�c�G?<�я���>�R���ɏ����
˳W�e�]aS�x}��]q���1ꐚF��Z��M3L�^۩����A�}�5W��� b�5�2�m�*͓�^���"(�"��7�q�1���`�{k/P~��Ū�F�K+w|�$P���<Y�-����;a�k���w��\�*!�t�o	�{�+s	����{���Bjb�5��p��Yd��_��F�(����m<BV�'���)��{C��mn�����;>د��a'����6�:�t�����^ӫ[Y龑��ѭ�찍R��F������E�t��4[2���y���6]�p������k ?�G�s���Nd�܈�m�ڏ8�������t}{�Y�T����ST��vB�&q�u��
Kt�a��T����'v�; "�Mj�0������-��|,�i��ʆg]�6��hs�C�~ST�c!�
c���J�(���OS�Ϳ{Q��7���Ъ��h�J�(��DY!������� �"�Xn<����c9��+�ЇG���D��0��M�
Э�fh���m&�;��̍��&tK,��,+?�ߛ!LF1M/��!a�������?�%(V8���-"�CW��g
G��ޖE��	�ds�v����"Z
d�����d��4�6[����
*8qU�s9<�Ĵ�`�����~{v>�]��4W��R���c��G����JjJ{|f[ ��so-��z����ԯ~d��\��������&�|~�4���lb.(�MTn�������
�u݋4d.]��vC_�5(3iy0�j	����(�l�d�~�i�_�
�;����S�W#�DvY�몵����Y��(f�"kѮ���7�Ն�}�������q:�B��\䈔��}`f/U7#�L����:o .2�G���^0PIG�@h�1��Ͼw�ky]E�꫺TԻ#�S���� �t�Ufb���f��J�)wC�f�.re�@ ӏ���#��N������Ftߥ��;��%�w�匫	-qe��).�y\Du�l��P#���H��?���
���o��i�^���m���j/�;[/�#�"��/k�< 3��l�"�
��)� g�ke���3��,0���E<z5�B�Cy�8�*"=EO�N�yl��xΈZ�z�~��3)��/��^�5�Q�Bt�qnz�� ,��&�0� ϕv��r���O���r��Ś\��|��0��AҨ6�ʲ�z"S���3���Cz�nqգ.��P��{��2����o�(�qgI�󪸤���!\�r� ]�~b�
1�*[���xZ�1U�ol��sT3,	̛��r�xu�[P�dP�5���i�u��'��q8zư����PHd�,ה�bJ��r��URIfÀn��|n�C�L�K'�����1��"!͏�p<�l�V!�.�؏�aD�*?��3��ί���C��r�Hx��U��V<��p�
�+J�"�1&�qr���45���-Tm�X�C7���8����A�j�Ǒ��3>I�h`PSG�D��)��t�=�>I��K��$lI����y5�n�������Th�/�C��Nڔ5�\�Lΐ�b<4��ј��? F{w��2���
ŧrO��N�$�-���'��{~T7���p��F��?�vP~��W�@��&^�E�O�@��Ȃ>7؎7��]C��92]G���I���ˎl"�ă�*��?-f�)Rr1?�����S㢻��cJ+$��@ B:������˜s4Y���sF�zm3{v�I��S�h�+���ܯ�as���΀��ӕ�
+�hu��9;DK��Et_�4�.��`m�r�e�`�<~I?L$7ᾚ�}�f#��%��pY�5̜�%r��V���WK��Y2��J�4f�Ch/?O!�^�ց�#�#&oQ�@��6mRkeo���Y8c��[ɮ�Ň��*�}���ޕ����|���?��poQ��W��%f~�2mk����]����aL�Ϋ(&�o���L�Ѻ-��z_��fh�m�w�P3'Q}gw������P!��7D� �8�{@vb����n`5.��k�E����������:8m��/����>�<(���!������&��817K#ԑPs��(OA�9���Q<PU���墝�����k�����X�Sa��:!�Z�a��u%Z8�{�_Y;A��~��2K!�̘��-M2:������{�k��w���B]\���{r�5-M%�6d�?uS�T�FV�M0a� ?�'[\W��é�q�j��gY����������ǅ�4��Ap94���FѪ^K�Y��ŻK���H*�N&�Bd-AcM�X� �j���[�;����$Z������F��/�t�l+��o��+~�����"��'K!�K����G��FZ,'��r�%`h١_4�;\���R?O� @aCm�¿�_s"�ԭ��A=��	�J���	��<��(��zW�W_U�	_�c������xF�q���dw�. �/���uE��v�Ws,���e�Y?pE�-��,(�ap��u�����NC��6C\G�+�:wu��yעi*2�~>���,���KFG.%<X�Y����+�E�^�9�V
��w-����?�ٮt$$�*�ef��	��]��۳kҢ�º�y	��'ME�����>ڬ�ߘ����:Y��0��L���D+K9q�9�:�Qb�a�j ی����3QKڨ(�v|�E��{�����Ѷ�D��z�g��q���!����+�9zN�/�= �('�o���\jN�<�\�С��.-ͽ*˥���^�g4Q�G��w֧Ix������^��$3A�g�/3��$~W��p2�������>���Kk�$!L(Hʈ����:�f ��Ӆ<�6ĲpM�ZՏf��^��齆@N`6�<�%ZEF����F.-SK�!Y�����6=�md|H�V���RU.B]��C�O�4��݈:����k�� �;M�<��ʃ���Q��\a�l����f�/�X��5Fn�#����1C�V&�nY����^6X��;N�����~$�YW��H9�|�w_�Y+�sQ�}�"��ܝ�vi�Qls+|T��d����G.���c��.uk�m����(��Sc/���C^XY�Fa�^�pO~W�b�Y�{�|J�\!��KI�$M��$�����F�Βlp�fBy��;��y%zjj�&��c-��	->���f��x�P�Ƴb�1��$�3�q� ;������xe
�7�P�ciO��׫b�I����S�H�O��|�ةi@��FUhkqO��"bE0�:Cr���%l���r	���%�Q�}`}��82C�]Z������Kj����Q9{�Kx�v��^KSln��]|R����c��_�#8A�������� �ݳ(��6��3즊-�W��+5W1;xMtY��VC&�M�'m�[�"�$�����M��d
�Kt���{ˤy�Sw���2��.�w]&t1ha*$�u2�O�:$+�#xۜ�;���_	�o_˷�`P�n��jV�/o����~��/�puT�
�D1GC�`~ܞ�hM^�V�P$~�)�0^'�<�ќ�PQ?�E3����V��]ds.:���L���,��3�՜3�����y�ƯW�B��Wʀ�\&�c����ۋFy�~� �s�Y����j	�2��W+lQX2:g�f��:�S5�^<1W��d�f9+/��fo+���Y�eRB=6l�<�s[��ܤ��œ}��U��'q�l{G�B7��r��5�A�/�f���{�-�?��=�R���v�-��F�Rd�e��z�������O͎��K��t�\{�I%4ۆ�7��o˔?]`�W��p�d��C�%�$f2E����A�	K�@ܪ�e�\ļ�ɖ����S�!�X���gII��c��{���������ܩu���^*̞A}�m�����r�`/�J��xBnR(dH_��3�)I~뗿!p����jU�p��I㞬D��_�	n�s~}�� �|����*.���@~
Qμ�jI�TH��dޒ��\$�A��I<7f^Z����j�EJ�ӌЬ�q܍ Su��S=�k|�J�g�쯺JȒY�ӱo�estϡq�F�GX��0����mL"�/ IA��Ĝ�{�����8w�w��s�C.o�c5dT���gQb-���ƂP�����#Zٞa�F%�^�20t=1��1~�m�lg{$�M�c܊�ۘ�B'l|��{d=���2���*(�� ����t��ȡr�-���"K�'�4��,��	\1��1�zYE�t�~��v�#7 f�.�0M��b%v�hd��ǀ�m�^�N(]@�����=�}D�}��h�.`��q�{����ϱB��E�i��NOW<:�Y������l�c�HcQ_��Rx�m.��S���7�����$Z@3����*!.�WH����^�����Ɖ���1O�Vj��s�ү�Z��R��/C���*���cM���Y���_����;��M�nbSHc~�"�72��um���1���x�!,����(�v����CQ�/�9���A��t��������/�2ٕ����K�N�3���_wxrP���Ǖ��RP�n^qK��,����V8n`[���h�8� M �l�v�*Dq2�T]��=�ƕ�|������dAME7kы�i��������(��ǝ���AFH��j�'�h���p�
,���"�[��r��W	N�q#��(6S��h%��v��'�����6pw�)����zx���sg؈�E���Rڊq�vj�l��1��C��fA�����L4�܃����9C��9���	�`�f��8�������:�}u�\2�,�X3%��)R�Gy�A��g�6����T	]5��t�`�K���u��)P��4M��k��C�D|�
?��g�o��W�Z����AQǅ�L�X���E!/��&Ou�)�9�i��I׿�X>��МX/\�9��!,P&_T_i�B�`�]�\�>g��?i������βBjɏ�Arhz�h����>�������2.K85�`6��T*�y�	�U8���S��q��{ ��e
b���R&���������S�]8�6^�������9�DCi�Y�qQ�� ��~"�zC7ؾ���4�J"�_��j���e�D�"̢��p	���i��H� �23yb�S/f��[˔�Qb���A���w��8�C�*���n�� s����:T+$}�5A����O��t;,�-�fC�7��5��>����ط����o��3.�/��E*SgȄ��ļ�h��T�g�N�!��G��٪�Լ��*��)!Fu?����m@���^HcnhC��5a��('��U6[�t'�*��I$�j��i�Z��;�$���G�\v�~��QAB��~@#���[�ud���ə��*j
n�­�1�{���_S)b�������@A2�78��7��K��)��*�	ʐ�G��BUޙj;�Z>C׻�q\hJ�|��u/|�I�U��� N��p��/9�k��,�#%����>ʹ�Ӎ0�*Ay�����$�<^R���DB�u��U��S�k�j�����2,w���F���~z�\y��#?�8|�4L�ϐ+��M1����%��Nڰ$�0���]�bR$!Xש��öipe\�C�!�j)���5�0��=���0�3�8�)�=��:�֊L)�m���^t�T��1�ހ�p2"Ѭ�n�U'ZC��0;?P�B%��P��s*�J��`��B�`�w�m-yBy�H5��+��ʕpҰKSZ���T&�D�?'�x�:H�~�
Q���7�f��O6-;����,��y�������:)/����`����<B�\̨J�4���	VI��50��ѱ�3����q4da�!
�W�\��׉�z�dk|�?r��^o-,���p?��Nl������
�x�B��/$��9}f�Sܦ`Mo�Ր�S#3}Hޭ4=���Вr�c�'{M���J���y����]"˂4cxb���mpm�Vq�.v���2�z���n+������%�*�Ƹ×�7]�?��Oa�X]��roY�r� }�hJ:�k�'tO"�E�E4w7 ����ŃUG�����
]�Z��F���}k�˷hb`Ɠ�A�R�y��xU��)I�o"P2�=������N�ƃ<6���'~*��۸s�-/k`b���(q�����D<���1Z��>��Ě�1�g�ʐ��@�E%�L$�O��a���l�+7X-F��zwǄh"25�����-?���r#z_X�r$ّ�޸�(1��5�U�ũ��Kc�}W���}yI��z������:ND�����?� ?<�\e��|}��r�\Xl��.jA�����v��iy���6���!L�Xf�K�������'�t�2�,��d�{���;^�xq�)G}�hP�tR�44iIn�QQ���Π*8S/���A�w�#��7���+�h�K6���ʌ5��ٕ��Mo���CHO��<��]�y��t��B�d<�g.X�<�C�Ţa6?�@�ө��"�� ���R�C���񺐊�q@Yᛞc��؄=("?E9/���D0!/Q�RQ+���ȫݔ��%v���W��@�[RP�daO��S����v�	�����CJ*L�2��J�Ԫ��1��u�!�t�<��g;A��S���<'����>)vaXŸ	�hPV4��<F��l;���AR>�JcR"��>�ތ"<� ;��z=V�(0:�Q�e&����SO��P����F�t�?�*WW��S�~��5�}Xr�`R1�H��KrV1��8�9��\��I
	�&�VC[7�s�f�)��S�]��AX�8TH��c�r�s��o�gX5�?��Ju�-���H�5�N��C7�5 ���?�l;�݀į��X+�⤘4گ���*�un�E��dl�G�ƪ-��RM}<mx��w���v��Y���CM�F�;_-!>��K�Q�����?�	��⛔�.�le�*8%xz�]���1����C_��SEk
�o�F�~k�<|hC��c��E��뙋}������ҩ6ӌ��]����<��CCS���[�e�E-�9�*�`�Ģ��U�VT%��"&�װ�>�Y��(_R��z���h0�&�o���+r,|�R�u���m#�����=�]2i�"N���y�O\��f�S���ӇV��{+�z#���{�ѼQm�nO1"��um��
���V�q.
�]���E�8�6 ��W������] pZ�Q{�ـ��13�ۏ�o�V�at3g�aD�,p���3x�O��>�(>��
A-������
���2����@�mg��Lx�I����u����Ѝ��pKI��/I�+�����/�0v��Q�_�L4؁6k���B���7�$U�rߔ���]g~�����Oi�����ZtWƹ52f�/|Ͽ/O�����
Eœ0��M�\QP��SY�N�$ɤɽ;�m3�?�6��z�x7��� ��z�U=�*j��
z�=��W'�B���a�s2�p1�8�P��AYo��;8���{�<�a��:�F' G�\`�S8&���ӵ�)�L���M���Y�Pur���m��̳%�k|a]�N�ݣ�LR����]��O��,�e�e�@���P9�;xI�{�q�8pK��1���LNImS�X�yDc���M,��7�3����e�i~���k6�>�揋k����7Z���쇾���h��%�	R���bOn����9�*W���|�D�Z4|�XN��G�~<4��)�tiZT�؆+[F���4���`����~�?sB�m�i�֝0x��7?ke1U(��쌄Ԫ����q��aL���:�ْ���Ƿ��؉�����$q��<p�W�S�xK�4�F�n���J�K_Y!O#h[��u�L�C]Zg�ة�o܍��0*�iZ���ۍ<�J�������I�iF-���l\ڶi�������A���0 h�q�YF�|��ZREu��֚^ �e)pMp���}f��we�G�5�S�������5!c@s��\u���y=��aoU��2_�~ƣ	���K^�� UH������_W��܄�#�K�<?�?p��d�rB�N2��K@����,���}q8'$���Ȑ�2��j��EJة��&�R��νس��AlC�8mu�o�u���q�
4�B��!�0��u`��I�&���M�$�����p�#T��M�Q�H�Am� �����5 ���+���>�lB�MFj�����^��P�w<���@^�!������'X���Uj�����D2�Ǯy�Y�[n[-�r��-;���
֞	�B���3��*�t�-��K��A�V�(X,=��b^���{F��Ϸc��7X+M��q7q�r��+Kj鶚Z0��M���]�M�.:�9��g����0I�$�%��<��u��\��4b ���-��$$������.���x�~^*wp�S��j4Qqxv8Z�5�������œ�'��~Q�o�3��ECx!��ѧ��Z?��oٺ�|).�o�Ǟ6H�T�]$��"
�=)�~ް���"�۟�[H�מym�l�� |Ϙ�@i���/���ߟ�]� 8�K�eL�v%/�J��ռ�^�\�ݠ�A��!�ͳ��HCqO:���@L�6�o�ǃ��<��G�A��}�s�q�o��LC���X�K^�P��'k~�(��_E*L�ұ��5M
��ͻx��Y��L�XyE-e;F^No�rDF��^0o�WUl2}�虙"�^�HE��y��ЂL���ޣ��Z��P�,٥�l���?������S�pۤ�"�C��6B�mI����ce�eT��!���N�&��nJ�}A��v�U|������v�c�k5P�
�r�Dߟ7���p��<j���~�xr����.Cu΅�Ռ|,-&^)u��P�\��%���	�?��cƐ�(�-t�=!�ך��9ˬ��H�wEd��܏d�D%�a1���W*k���[c�<ʬ,�l�xr��p�v֒>���w�I�$C�a�~m�8Vr���*����-)�ފIZJ=iu�M/���B�$�b���k��H���Ì��t��TZ�i��,��=�8����;��Ȱh�q���_�r|�8Q���~5����=����ttQ�7��q1�ot�ء�/'D�x����O��b�  �"����:������1Μ@���<��P�P��M�:0N�N¤���L�Z�|B`�p�lA���rVrd�"�g�paK ~�A�e��g)�oƵ�*��L�j�*׻l��ڏ�9$pA��}*�i2�\rm-�𕋪K�����/�Ӝb���T���*�M��zi(��.fx�/ԕ^�1���ě�T 󟠸�`��"�ۯ̥P�A���iqK>;pc�4��iS��3��K�@��0]�����o��׬��J�`ƛ�a�ڼ㵪��?�dZ��X��w=3����b���ō�\9���S�Ʃ�:�d�w�J��z����x�+E�3u��O\	�m�w-Bj$�hUvj�U���x��g�ϱ�
39�;��e3�O�:�O�U��sV�[Wu!��U���ղ�F�n���é�T��2���%�b �0v����ꬊ�-����b�9k�"y�eVP�K��߰e-�m��mMf���kz4F�j�0Hi󻋬�?�(K��,%KE�^ΆJ�c9"�6�R�z���Xgg���v�D�pG+}�6����|��^�����>6 ���A�k_>�}wm[W�Ô�R�E��*���w`Ns�[�ɉ�'�j'��Z�E�F�N��:G�lc�4c���jb�h3�cK`���?2"X�:簲����e~�L�1����%d���Na���H�e�x��vJ�C��m;���ځ����aj�{Dtl��o��*���S��u�M��q��jbX��9(�r�xG� ���t=T�
�a���ժ�Vf��Ԓ5�::��Zo,U��&凝~���2�����We�hٟ}j�Gh����O�1�Wӡ��;�����s��P�2������EpX���� �����|��Sh�W�G���t6T%����p)lI�k��EN�-U�ym�E�3&`A-�.q��=n�!��f~��ԯ_��/ѻL��9&85K�ר�X���_v*a'��7��~�!�E�N�ŝ!��u��|PT�&/�oO�
�0��{q"U���\�ߊ5��4�Z�n�Z/Y;⯃!����w>��2�r�K�|Z9�1��  ��ŏ>�<$q�r���t�U k^��){r��aP��*t�(��F�T�G��%�E�S�Dς��Ґ����PF}�sj��<��6��}�X;��WJ��Ʈ�PK��:��w���Y��B�f|6_�?�u'�(M��H�Z�cV,Lj��B<5 ��=�&Sx�ʡt@T�2��`��/iiB���>�EC���T�m&t�/����{?��5�Ne}��%��9��[Pc�A����j�}�dpΛ�8:�R���;٬$1)���3��y+5{KPA�!��eJ��D�mG���!#��ژ��D����߸��
�\o"z���,�ؼٟ�ة{�����+���SΏ��>3���屬$�;"�g_qPi%L�>��?�BD�N��ު��1��g%��9(�U?�[#�op�HG��Bv�:���!����]���Di{��]g��Rmj%}6�<30����<�/3����@�Y��ƌ��k�B�9	�j�r��V��X�!)V�Z�~YM��������J�X�~p!�� �?���g�>��%����PP�̀�F��.f	�);�F�s��#ç�=���B*�qr>G;^Dvm=��F����p��Y��E�$�A�c��.+�uW��@�o;¾iw�[���&��/M���)V�� �kp��1v|�Њ�] ���O�G���� �8�]�	�9�����R�+���9��P��*Y� A49VNZg9;�o�	5����:��N�Lk����B���3�F�N�s��-f��p�2�Mhא�3�e�Аi�q[�pM�ɛ�j�r�19+��$�C��&Q��@d-�Ĕ6���%�o�]t}R��޺׺�Τ*�(AMuQJD���ν�Fl��bI;�4�T|�uv���	�b8gh�LP�S�|�4,ED��"^�������8����J��X��d����9Ʌ�gM��,:7����=���YhĘ�h�/��i����rE����.���_��b�$f�3H�Dp�]a�&A�S�ǻ�t:���e����
:�x{i�k��c��뜟7�@����$�;�?�4�y)^�!9��}�SVFu��,��F��3~ҿ���h���h�]�shB���^�P�Q�CL��W�"P8�Da9@;h��W����F���ic'5�zW+��#H��J)�<eĸ��**�3���}CFz��2��$4L���W�T�G�F���$��L��Z/h�v|�v�C kȇ����?��&�rmNa �P��$qe���.�1U��ߔ��"~n����z/>n�ϯ=�>[K��4B.����ǀ
�!5�|y��\6'g�!ZD��}���  �A~i���z��S��k(%&�d߰�fY�L��+.�.�Ym#���tz^H��A�Rh��n͛�k��;��)D�Ѽ�� Q��: Z��E�u6�q)�3�viJWa<�����5��>�m3j2�:����exob8�t����e?�/�'|�YI�x�bْΕ~;D��x6};K2L�*3��MOo�܌G�{G��G���T�N��s3��]�)D��n���ޑ�����ҏ]�To���ij�W����VG����5fN�,�Vpx��CWO�|��4�q��;Q��U�In60�wBLl t�#:j�����N#]���UaOR��H�9��-���c$|�m�e}YoSE�S��P���3ٱ�l"�\K��.~���A���8�B����#
$�PK
��<���5��.����
��<�n
u	���[���G�7�{Vp!M��
��V�-�j?���2#�+�9�;I� ��d�{B�X�ű!�kU���]�j�2�w���S�KwT� "�(�s�O���HZ �̥pA��=���;�1�.q �p`s��(/��0��ư�/�3���ѸDXo4��dz�f~���3e����#�录�oצ᳠`�����`�dڇ�{� Gّ
1��\L�t%L�A�zk�0��@6.�Q��,���Y`�/�^0g:�8U��Z�[�=��q�I���{�ބ������3��&U���eUS��J���z���z�/�L�O����L�|[riې���B�&�\�ƞ�{�P`��v�8!��Nu�L�;\����hN�ǎ.����$	~�g�栈���Ҹ�/�ﶧ�ll�[���<�X�Y%^d��M-��8r��7�}ʋ�\���B^�������-_UB�!"l�E���|�\����8�Z�Qp��&�~�l�ߧLN���e�ŷ)���Wչ)��i%y��V�D�:|�޺�D�J�c�v����[8�993&�d��Jƨ1݈bM�q�ݮ8�Y��촄���i�?�c�^�k<n�h��yD20�|Hu�K�U�p�@�(�r�$���THu��+*^}�o�q�ԩ�@�v�F}� �%)QbtGQ(sR�d!ί�/ D�Z�k�Oo%���9ɶ��6g�z�L<P�5C�s��Xfu�Τ⎃;'�z2U=|.�n.V��4&o�{�?�B�ᶂ�w���ۇl�H�{�t�Bʗ=�Z�(��t�i=n�廏$��[�
���C�N�d;�?�c)FR�<�ec�R�"VH-�̸	��s�
7ͳ���T��;�y���L�6��F":��X"��/�a5"�R��lSd�+�P���I2� ���r���29��,v&����v �3n������D�ua�T��\	����܍��^��	�H5�m��5��w(=���<V��0�p���+��bh�X���y§�`g)if��ܢ���bpQL��S��șג?��3�W��I<J[aWqK��qY8��d��{BR]����0���0"����p��׌���:<�I�>�D����1�N:d/�H�B��~���>M��h7�h�&��m��e�L9F)�FӜe��o���J�|+��[��rd{�+�g��1n6̆�HǛi��
$Ǌ[X�Z�9��f�A�W�;�����#�-���B���Qx7���o&�O�>�jF�o2���?�\|���r������4�������)���S32/�Ī(�vY�*�	؈��NԞ�S�o��{�촋���������F�o�(�<�M��ʈ	��Z[yo�3d+��j(��zU'W�|䗛�������&���D��[��Y7v�����J��Ϗޣ@����~M��C]���+q譡䭴�����o�v�.5X鮽 |�6'� ��ʱMVқ�
Zm:>��CDJP �.W��P;@4����i�]����E��[�v��O1drgo�Ο��Ѽ?��p��4��QЏp�����<_�$a�%�|���%+e� w�ᇩu��6��-�b����U$aV0A'��f�H��[�.���E���qz�uZW4\TR�`=��@�}"~�"g��g<�`���Ddm��/�DgC�g�(��U�=�;�e�>���U'̖�!��,�4��M-H K� j������3��Q�q1����ۧ���_���NQ�XA�:��d�d�A�$GF o[�D!��X��at��#��O����l��"��f;|����쬯q'��/
b%�zY�2���:�]ҠŦ��\�z_�-�;������0q�2��8">0����G�*�7��|����# �.��$�5x+�f��C�C��p
�"H����q&�"Y���x�y��{����F�D:�gD�6.����J9���@��o���,>��nqFt���X6�TlK���ﭲ�����;4���a`J7;sku7��{�X��r�F�~.iy5?�D�<m<����V-+'fu���F�hU�mV����eF` ƽ� ���s����aX�^X�Ԛu�k�ɫ+�A,��=�Z��f{E�9�!��=uk��A��K]��O�I&I��6�n�nG��,��s!G�s�0��tIc�Q�����������s����?E��M���Ā��k�#&��E-R�s���O#Z�o��T�����/���N Ё,�����(-H��b��\arGãi\�XN8��H�L-��f:�k��D;2b���lav/ �%a�I�8,��0M����;���݁��M
���իj/K���^l�������0b��y@Y�{�����`�?$^�Y��&_ddP������L��<~!��32�<�嵮�1�Z@k��8�������1��ZqS	�� ����ʤ^#�CY5�FܠA6Y�KTz+ڍ���f���2���}&�(�˞�>���h��SH�)G� ������q���c��O�A�g4"��c~"��+�M)���S�,Pt�i�Ƌ[�@n%�� ׆s�0(�'j^��wc�����JO�^� zS�d�C�	C���h�d}�q�1X�&b:���v�����ː�Z>���AYH��!�[_):��� ����5J�}�b!0l+H��BZ�z�r3-䒱��޽Ţ_a�ᜓ�[�tQ��?�[,�֕8hH�b��G��@$��i���Q�)�Uly~X4�j�h��Ѕ�)�zV�m�)̉@;!}�m�=��3`=�lü��t�J%GJ�d�H��/��.8��o��ܤ�z+�)�4�n�I�r!$���Y7� K�q*���<ۅ�I���T����H�K:UQU�R��T�:�@�R0�رp�C\-b�<��D�gWR5+-P�de��H�3�*���s	X�������
㛍e�y��a���G�ɻ����B���Ш8�ܚ�\�MF�}f��Q�.9�`4��֗:PP���m�c4����Ӑ�dJ�Dota(���U�ϰf��mi]�ޙ�IA��es�f���,�|�DDC!�Ʒdbv*�Y*[Du�{ �=�Ņ�c��� �����?�%%%�K�}��>)�F�6�����,�6/���ë�	��B
sk���K4�{�Y�o���W2���l�q�%����4��Ks��5	��0PW)�����;[F��T���g������T~^�E�a��ه0R�K�տ%�]�O��}��` B앶H��G���m�Lr�|��&���EM;&�F�5:h�/�,���B�Q&�Sjd���si|l�p�*\B��Z�{�{W��\6S�w���M͌�H�U�����Jas3����1��>�����]? ���=�wd�b��� �����F��3+9$9%�E����ڞ�=>|���5���NJ��\��x��o糂�SYu� 7��	�����q,(��.nl��4 gy<����r� S�9����J�?��۽�����+��V���Y)&F���� ��\NM`��!kIdJ:B	"Q�����!@�p?@�>#��u%fc����]6$yo�K�m�����	3��Zr��S
��������\��8ܒ��xf@�+a���i�o�r�M��B�.FG۷E��<�u�(x(,��5A�S�$�J��[m�Ց�z�1��鶉����}ARu�(j�䑿4���bKP�A7_��s�PDS��>��?8=G�tC9&	"��{k���\ʀ�7��j�"_p��;�4d� ��]�x���	�i.{!�$G��;�"�z�C�
����]��Tvݦ��c;b����h���j��D.��Y������W����H���!5��c_N�Ⱥ��=]�Go�MG����{e��{���E}N���.O�B�3h�=���&QW��������o�h&���C�\R.~��
-���	��E(d���Y�Xp_�-D�Y�g�5��N�4����9����+��:P@�9�-H���%�
�X��Z�i�.:����O�|�_�/���Q��j��۴i������9l����
�����3ּ������6L>�\�N�Nb�e-��h.��]A��qa�D�?L�O�y�/�@�gw���:5Fƕo����?5 i-��g�ʂ�����j�����Μ9s4M�!��;̾J�a�l�2�ofP�.�Y�̵������DVN���-�H���k9́�7{YW�,�O#��K��ȫ�T���#"��2�yS=)~��.n~g�ne�҂Nm�~�(�澁%:\+T��?����%�Z�'5t��#�b*��sF�M��XQ����$	�/�&�P�f� ��Xu�� A�Q�����'�a�!}6N\'��P��h�b��/șȞ����{]�ǚ��ݤ[PU4����r�Q���1���9����`���U�pl��$ق��#� �	6�:)HY��E��1�PN0�y�e2�YTZ��z����Wj�V�~��=/O's�A7�9�I�2�/n����q��B9�#aT* �89�u	��[���F�L�8��o���a�Z�Pa�KV�)�c3͂ 2���RU���GI�"�JQ�u�b���}ʻ���EeG8��Z��O|�D��\�<��sĘ.�[G���L�IGAK��������KpO�������.m0��|J��lf"E�ե�!���|	��!��L����Df�������+	Kh�4��8u����7�4��IT�B���z%Re���֠���f�T��﫹�.-��������` ߪ�EJC7)��o_��#sѦ��\��7��Wy�0��F���X��e�l��/�0�(��n��u:��I��r�/a0�Z�f�e�T��pcVU�DFJh�o�i�+Jy����*TD��񯨢�ԦUeD'�d�Ö *upn�zM�R�FG|�V�V�:(''!�3<'$`9�F�r��w4�	�34d2]�2B������u�c���j��R���ꗹ<U���=J��0}4�g.�	!�Ϳ��p,���q�Ɇ<�� uH��+��m�i��.p���k�2xP�;���$��KbZ�t|] eW�8�}��$b�Y����1M�J����)�-���Qr����ee�ڮ8g��O?whs��8`<[Y<�1Q�ro-� ��I�Q٣.�阰��CA,�P2�[�fD��Jt@T.@����@>
{ci^�p�D�u��4���d�3�h�v=y�f�(4טP����������(��⚊O;*R`�BExo�D�,C8����oAۗr*��p�54-�0�t��6����{J֠%0�z%̫�j�C9~l���/]\�G�����`8!gP�8���Fh]*�}!��5��@Z-����Ȯ5��S���3#1[�G�Z�Rw�]�=9���7�G��Aã�Dd?Im�ߑk=�}�1�q�^jP&F>�"!x�&|?��ޭ��W�1�Ј[�2�x�4��KaW/�]AI��QY]���F�Q�l=��
?ٗ���v)�s�r)ƌS�Yx/�����iVC[�3���́G�bVc<�	��F���R)�&�!ϟ�=���q�1x�l(l��6� ��K��!v���{���K��:���"�d�@��hF�)jle8[��S=����,��<<"K�N��o�B�+�Q�en,�r�3�:U��iz�� Ɂ�Ⱦ�O�$��OQpE�%g>}ʭʄ�h�>�d�H�ɼ��5�+;�`Q#�p�p�K[28}�6��e+���P~�Yh'����_��e�Ƌ4����,a������h�VM���/���".�C��@r#r�Qo�K��Wb�=�Z$��~��nlԖv;�0��l��H ��Ƣ:rJl4�@��抴EZ�p�C�����$��^KFt��=�GKfW�X�P�꼠�?���'����m�C�����Ȯջ��8P?�"lUc��a�UxA��g(�ضOjG�Lᓘ�1�(^�E��[�t�rt��WY'�������Km�c��Fn���)g�D:8E2��ޭy�frc.�h�G8³�m��5�뚐Q�/�Y�L9f�׊"��'�j΅YJ�S#�9���$�:8y<*�yk����]�G���ǿ�,}�no��u=��<��9��;���y-�vZ����I�?	��Ǒ�{P��/������SPxh@A"*럃��a�z�\�ߪ��0����_�י~���!0c�� 2l9�քS�(d�'gS����}<0�c�`��#�F�*�Ȇ����H�R�����쟤.�0f�F�u�U��;�:�]I��
'�`;8��2US-�$�(Vf)6�)J��0���y��N@F��9Q�06��g�iVj�2��}�|Gƒ|�ovd,�hN���$�����FA�شu'-.r)��9M*�����"��[��J��Q��Z;B�O� ���������'PO�C���x�	���U��X�S�{��"&��AH<���X�L�te�b|Zs�
Ɉr<*@��,^�Z����Yo,���d��ÄJM��#:�� �_G����Utg�����ꥹS?a�[�;9\f���k��ɠ�1<�Ϥ�:����f*)�֥G�Y���h�CV�iI 2N.&Qzq_�G�F,t��Ai8;��뚕����""�Q�!�D����� ���<�ų� N�}{���D� �R���]<��徂ӳG��[R�>석�:��6t"���"T��Hpt�����lu�E����<t��de��\��)14�7�W9;��� �pf�ײ�3�GLA&�eA2�:���M�߃[g��'ܪ�l�U���S���gI��B����p�V��Ǔ 8Ky{8�'6��Ff�8va����x���v�/.d����5����y	�{���z��_�n0�w���m7N�=T5X��a'��k��Z��/Qإ���FD����9k��ȝ9��IO�*�l�T<�F�i�s�&���󅯥��;-~ڈ�&1=m����DM G�6�o�?�T����U�1�� �Ap����״�0֮=5�M���x�S�����>c��X�?����,f�kKZ�&b�G���Ц{>����l��dm�]�ڿS�7��M��܅����L���,�#K�JeL�!-��� ��܍����g���/'Uuө��xE�Bh�e�l���Z�����V���A�D:\��(:4�KݶV�r�@Td�E�6��Cnx/�,���2B�t辅t\4W�%��P"�ț3L�.������^���͋'	Ê���������M3<���j(BmXuq2
���ĸ�.WU]�d�+����hn;.�vE�jQ��B�x�𒀩�戝�8J�ٚ���7�9��tE}�4�;�Ħ��ւA�s�un��G^��z��v�b�H�$jY�4g�C����*t�������;#��8�Ĕ1ąLƷ�Y�́he���_گ|gr1���.�W=����:����*e���G�3�����R���C�`FˋKw"���y�TB��u��<^>oO���U��?8d{ܲ!ǁQ��I��?S�����gCu�o�R�7[F�*Ɍ��A��ߔz�9]�1� �ZA���K��X�����O��t�YpϢ�q }�ɪ7�� ��`��]�5����$O]�9��%"eZ��8b�|M���{%��^�G�Ǌ����0l��`�eՒ��D��j�Fe�G�9ZYT>zu�m����̢V�9����G�T�o�EJH���O��0��&p�V4b3VpYĥ�9-
�J�}�:4'us�3q%�5!uO�����@ghBp궪O�c�I�E�8�&R}*4����p�_%��}�'}��(;���7�?����B�:���� 'z�d�v�o���biXG�Z�Bdf�x�~	p��(t���U�5���w��*�}�8�o�������Ԓ��;�]M/��}�#�~�H�râ���n-u��^�o,�x�a�f);N�G���lG��q�l7w��%��C���"?BzɪaZ�g]�s���
ӏ�ˤ�zX�?#�GKG*#�W�V�	nZ�3�����G�;��/ʨ�[�#+���{���翐�����Ҕ}��ֻ�Hl�{���߾ࣽƵ������zβz'��(�hջ��Hߦc Ĕ��oe���"��\x�8�Y��Nw�q_s�y܉����7|{��@d���11^�t��j�P��Jw0Ѳ�-��F�ۍ�f�$�����(N �j[7Ro�C��)��1���3�d����K}ޔi��D��Ԫ6g��C���\g���l�W���G_F�q���L�s�(ą�\�}��C��i���v��+�L�V��m��~x����O��~Ɠ��t��j� !J�rt]Z�T�YZ�X�2��\����ƾ��4\�{��"���v;Dxx��ei��q�F}CM3�ɉ��c�*�!�%vI�j ���@�8H�����+�	a������_�^)�`%#rgR4.q	�����ڽ s�G�TyX�I���G=L?� �2��A�M���E]$�wH1R\�C3������A �yY.��"���F�TW�k!�~1gm�-��F�9|�E-�dM?�ms�m>Ħ�Y�0��1�����b��u��>=̆�k3���E�����P���{	�9)���'4J��b�A4� ��T0��3̐�� �p���ZI���l9�|�#��ԴC>@�'He�J���`�.q^+�d���3bti5��G�������j�_N���t��r�-}��zw�u���qp�JF��=��h
��W`g[WK��zX\#n�F$���L}�����Qw�c<~��������T��"�#�+{��+4����St���[;���������~� ������!|[�Z���P<��`���:^�ՙ�u����`���Em��
�h�_�P�KU�F ��d�3��!�q?b�}7+����-�c�.t�����H�Z��)=ep��C�zŁY�c��=�<�Uݡ^�`��6��=�Vz��$d_��_�/�J2_����Ŧ����1�o�^�7SL��Bo~[�"D�#���2�IO��ա�5��M�p�,?����Ln׿�����*0�v��*a���L~��Ai��\��$K^�DC����=��C<
��I���	���%���X���}�3{�ߒ�x=��x�>#���ր&<�/���Wg�F�{�^O�h\�8�)�����Rp�~��uNԪ:M)��F�i$��u�p�@v3!��r���o�L_�,��ĢǙ�3ʭ =�rv[IcJb��+�����u�&�.�;�`x�X�e��aE�]�����֍^��༖U�̞�!)��<y��:����dY_-E$�W���Ŧ4��Vb	)�Mi'�R8���>�8��&�3j<L��0K��
hbw�r�c�9�a���\#E�|��DT
dO��[SV������W��O�Wb��y56�3Yא7�K��E��׭�ik��9��&FuH *80x_*�|_�Q�Y���Vb-������!��Y�HNo?$,:L[}�.�V7',E	�E�N�:���K��|�0�g(���̕a�6~J	l?=��hu<�j��4��ȿU�5���&UQ�����j���8��d<1�+���)D����T��g�!v��~�G�X5�ײ����8�T�;�@{��E�7}��Q���4��>�m�O0�x&�[SǴ��,��?��*�*�!�	���Ca�!��[;�U����)�`J8�H�;���$��u�Dh��❧[�`�tL�;���f����hrX�G��'Ϳ�uC:h�p'���)c�!�<���B�U�ż[�П��.��$��LƏ�BA{@r<"�[/��e�kF���[;�M�����j�O/n�ViU�c1s�L�}6�S�}�-�i0�>Q1��v����AɹW���:ӊ��65CL�8�Y��-1����Ǐ�4�����=I:�$�?z5�X$�5������5�y�%��8j\��H�Y�q^���"�I��j"��>�?����	���uT�
���|� fԝ����@����mZǴ�fR%��j����x
�� ?T̙��l���8�>J#������0`�]�" �xL�1b��{�'�Z���}τ:��噋|�+]<�e�q�����Z.�Y���_9M4P��-0�D��t9�ڌ�Ԥ�0/�$]κꗞ~O���S!�N�ʈl�M1*.��-�>ڻB	U�V*�[~��,�?3�΢<ĩ�!v��/�֒����f�f�IB��KwvA������z����.�J���W�Nu��Ο67NKZO�%�k�*���A� L�VX�y��D	��ATh��7��)�\
S�7���!�¨C�l�-(Za��%� �R�Hd�Wc�8�&�~5*�9�[	#kR�z��H��Q�����gu}�:{�A�"�<!I+R��	�Ҟ����*v~�5B�_��_8�JB�B�	���A�w�20��E�vY� 	}��S ���>4�`1�Áv�y��𤳼�g���F�U�lz�e} '�(��BVA��-�Dn���I�Z�Ms���V5�B� �s��5�Qk��ŷ�m�����K�I���&N������9��`Mlv0u�_�7�B[�G3!��Io���:H���x��"��/͖E��������P�mZ���^��1�`QזG��_��C�-%[��uA�)MK]F;֫w����0mz����6�_{�qw�ΦXDoZ�b��Ν;䠴4���]���(:�+�"N��m�	�P�w�G�J������L��q#cC�u(37��~u�j(����S����@Ë|&�~��'��v���u5�<7�s�)�;)��At���b�A�ڶGW+�Jp�D�&��HgOX�����7���_3%BFOexh��b���V3��o��9U� �q݋�^p5;��F}	�����|�a-Ry���e�f������P��J����t@윗����GK6L��)���=��Ds�0s%	/��P���/}��Y�GO t��=Jg.�I/��)1n���WϙD�i�Y���a2^���I��[����Nl���{��3Sn}�M�eQ�?Xe�Ү�[#~��LB�*	/�$�,��� @�1N�Ɲҷ�R������k ��l{IN���J*;����DhS��e���������i��oO�\C��͟\[�<���<mR2�a�b���&9����f��ЌbB���%��e���*N������T�����ZL��XL�9��ʓ��9GS�0H;�#��@�G���}��*�wT�
��!('tYv�i�k��YI����T�ڸF�=��_��,fm
�T!����.[��+JF|lǰ�i���R2�CWO��B�j��~�[W���t��%��(�.��3��s���K_�4t��I�|���� �PE�o��޶��P}��qy9^�*��ݹh��^��6�V�r��}�jl�IS6ao��?/2���"=="�}���"hǦ�6���
�8�H5���`��dD긤dر��Ӹ���V��7��<Է��9�$��"���r�M��:}x@6M�����4|#�".��ӽA�dI���M3A��#�}f�E� 	W�ؼ��e�ܭ����N:;�ҝs�[�Jh�$u��/�Yǧ=�g
�K�����)?�Q;톖��B"�z,��W}�[��w���<WzD����Ԫ���ؼ*㡔�X����j����1��u�~t8��I���5����L���Y�L>J���/��Ѻ`��=�8i7S��[���{Ls�D"V���Zb��MjE*���FS�>�#���8�cA,c]�օm�7����?���\i��������W�$�iy=y_��4=a��ߞ�'C�j�q��0�k¥�(t�mb,�E����]��Q�M�O�)�l�>5H' ���`�i��'�̝�z]y|�<���CO@<o<��r���`�Y�,��C�q�h��r_���v
��m F��ʃm	SsQPOk��inK�����o�f4΄�H�H�!E����ZņX6����=۱dT�=�%��S僲Ș�{e���X7�D2���P,�*W��]�%��>��`Y$�?֮&�%;�����#��w��K0�)��m{���
��
+���Ky������u$^['�*̀��b�NIA�Q���V�1U�n�O��޿�O���ɰ�"J�{��g�Ǧ;[0
N�1~�6��~�ⴣ�� �Aܠ��ϙ���Y��m�Nh݃ �!�O7gՍ>i��������/t�ү$����f?����},�P����v{��㟸�Ԉr�$�h�?JF���|�wa9�r�Uo����6:@������MeS�gz+6ul�$�r1��(�� �)��|P�� �_�]�d��c�˲tL4�:oiw�;��T�V*���|� 6Ȉ=���A_��c�a��s���M��N�*��bpҰo�P���?Mb�X~;[���@���Z;��������yjƥ��l�*�����E�y`���g,'�F�i��>�����b;��֩ ����cZ������W G��4(��Q#X������b9��N;� H�������hƤ�Vޚ�8�8<���0C�Z+��U5`��D��K��m�6pV�Aҩ�<�s��ӿi���#O��,���,��`u0Y��(������N%Yv��0�.�.��N��bL�h>�8݃�ϡ�i32$��T4W)9y~��?�1����No�kOS�S��;�ǽ��:��)HT�6�X�fAc��^Ӡg��p�9�M{U��qw¢�bLL��#�w|yl�gGD�,D��{�ر_Ӥ����I�7�y�ےt��w�硉��?�z�m���� b�ʆM��.*���g[b ���o�/�f#Q�l���xL�V��0���.<����7����e����n��H�����4y�X�g�!�v%��MkQ��Y+��Clo���4�
ʍj�3�n�X�i43�/&X/u\*BKHho�r��,"���aj%�S�Q%�V�&��"�d�1��6�e���ᬃJ���7\ɲ08t�.u��K.s�Rj�l�&�^vs�(�'��ªZ%wI!�5`<ܞ	��a���
�
6����ȟ<�N�.r{��d�-Z�&���ܘZ�'���mk�I�d�wzw븚Y���f}��4�?̷�]�m�%q��}��O�^�r\�:�E�:���$��K�Sٮv���*Qe�Ȃ���9��#�'Twz{��Q��	X� D{	aG�X7ӳe���-z=c��Q;�:��C�i-��n�(zF?�}4Sƿ¤��k��!�H�79���u�Lzt3*5�y�\����v��U�&/~U���ع�R1��E�A��:�2S+��/�c�vs�/��$zq �^��g��sE4Ok�w26�^��S�D�!W�~�VW}x\��|��&HX�y\7�<H�s�5Hlc8��s�Fvz�.,3;�����E�ߣy��s�G�r�J����}ˬ���#�H00��C��2i�ޙ�=�y������WhV��n'J�Y�B��yi@_��.��10�Y�L�d��g'�}�IR(�l�"�S����x�-EC}..�vF��� >�,}�$SX�����=ϡ��S�!������w�͘?|�p����
��K��d'�V-J���&�;1��z��i���?V����l"�J'�7����Y&���1N3?~�m���,�0��y�@F�f	����<#��|[q.���� C�@0�/��4�CD}D-�
�E��Վ�>�p8�����
���V6�{k��#tw�	8���נ�"I
1a1��q�y�iJ	'Ou�"���H�Mz����^�B	��pH�*��������N}$����Xs��Z��Uא�=[(g�a ��^Y��L[R�f�g�y;�Yn\�dz9U�;Tspó�� ���&n�#�n�X�o!%T�X�=s?V����i_�`�����H�� ��"Z�֨	]��H9�O�m#b}mG���
�>qk�}�*`�m�����%.i��*�M�o��y����p
z`�y��S?j�D���&��n���!�V��&�2�DK�3�#VZ?�) ��,��2�4F�t"�����M5����(��|��&(�;ˤ�7���S8��������P�zU���<�q��M���K�ؖ���h�N@�t�SӰ1��w��6��;����7�W����zR�T}��n���=t�����&�η]b�+�i���H��dhqu>�hi�zSyv��zlUZ�Px�&Q�~
��%+p7���sa]'��Z��Tt����{̀�Jm]��#*�p��i̸���&9}![IS�(?����jD� �W��] ��D���$��"��
���� 0����T���U;i�*���`����M��.�b=����� Yļ�B!Z��Ux
]���+ꩅn.�;�����|�+9Ve�W7It�깘p��� ��B��7>� ���������9�-�!a��ۖ�ix��P��^��9��� iR�;k'�՚>�"�D���O�j�H�����`?t18T>�b���(����C jv����KihD~%fG��C����	D�){���arcN�>R;��紭c��}��Tm���f�CF!Q�i�|d�,D���TY�<��כ����ǃ�'���a���y�yahb�������%W(��K
2T�mI���U�@ e3?�����#h]�'v���k�����R�z����M<�HG4a��s~u٦;W�d��^l���ٗv=��lW�2v�68�:��4�p8S!N
�������\Z4:@R�I32����X$B��gC� `?���\�s�K�k�r���at�
/���Q+OCĳ=�N��0�ʯ��� K+1\�]*�Ď��NS�/�v�C�̲���(�e���7�wnS��P즗�&~$}d�� �>�[��u��ҽ9�|��R��U{N�hB:?�T�)LI�7z _)
�J�'��m�'7(�FPܜ�7��^7�^���z�
�>�O�F�e7���{j��.�y)��7�M��O�g�1]�W˸:]��*8�\�9̬��q+պ��-�ĺ��쒼�� _�V�ea~�R�FE΃�������O<6��D9i#nJ�4��$+��0q+e���Z��/X?��K�"6?ӵ�.UJ��ǫ����E3x���r��RH��>xpUⲍ�p�����vchi=j{��g~����'������~?U�+4o�� P�%��4[W���M�=���o�>�{��<,�����>��l�et��"����]V�U�}N��5(c��*|vY��6�dS��x���6	Ț"��P��g�7+�1�@�]�P.�$(����}�,F�{��O�~�_���E:E^!Y��<�#/OY��M�q��9&s��e3Ke$Ip�ψ��F����<��k��Rm � 5}Z���m;�s�/"����,����%#�#yB�l=�ٺ��p��=�j��,��J�){ ,���җ?4s��Ko���c�Nv�z��j|���xj�+�|<���&W�Z�[h�C�����rq�P�wFp�K�Sd��Ԙ�H~�sx�.�&��B�sY:A�即v�4�V]2���D4J�"}����Іt��1͖�^�7��:/Y�N�Q)��x�&"�}e�[�:n�nu, #���&D+E���#k�=� U�4��Bz���R��[AT}����� �T0m���+.J	j�Q�r�3l0v>�:�[��������2������2��_�z)���ģv��[ڥ�4^͹֔_���Ŷɠ��m�m���3�c��Gm��G�J�	�_�!�լ�-i<~� S��H�sί�eeq6D.�*�	[D����I�e?�)�oTgWKègkFU����2�]]�-7���^4$euL)�Ĥ���6�N�c���L$��K����ɕ�ު�滮���ٸ"ѝ\��*)oc6�?�n���a���e"{O]
f%s3��I��),P~4�qp2�tЏ�a�s3��qW2fW
��կ#e�F��a��_T>�TS7���M�}��mC란;���U0.y�'����t�n�n��x��
��|E*�C2�]�e��TY�*�5+z���-�Y?��F�͘��6�M�TJrڅ~M�t�H��Pi��hȦ�W��5s���J~�&���� ��SGW�9��hr�Ɓs��*, ��u̝`3 �#Dȿf('�U����c�-�:.��M�9`π�=OӐ:]�l�M���K��b�����e��{7ږ���W[��]��?֤�W� 2`z���J�����#H�J��pg���^��]=L/�P�d�%��!C���TEw:��SPK���"���X�땧ŘZT8���f���q�%7N?쟠�߹����m-���h��#m�3v�
a6N�CD��9�i� ���۷��TT���kl갭�1[�����U���m�#�͞�f���#xgɃ��=�8��d?�A���͜�&˺�A�x�Ɯ�R]ŬO�0`h��X����1��T("=�o�|�օ�+8�x.5-W�����'l��;S0� "�����
��Y��.ݞ��h+���T���iFnz��~��9����2sJ�p�r��S��q�s7�_��{�c�ڀ��G��f����s)"O�-�(:�̸)�陥e�V��{5&������K��:�[0��/5�Ft���r���إM�%|���P�7l�*]S{�?	B�>$�S��;_�����4'�\��(��8��\T�3M6�_o���6K�)�Lp��n�=;�����+k���wB}���i3.��؀��c:^�P��:��p+��q�;.���O����n��U�>1�2����d��:���ؽŏ��s5W�T���"í��Zt�ĻB�&h�E�U�Tr3�.D�,�!�|�k��&3�t[���Dz@��?���@�Z�вg4
�T����o��A�Tvd����Oe�5�g��=�Ν�o٪?����q�-��9�*��c�;�@jT���lp&,5`����L�K�ҏv x�0� 7���V���7�zwik��]�N?Y�a}r�C��G�U5W�8��|K-�����Mzk����̿��᝽g� 1�Kk"/����v�)�QA��]���fTH��n#�^�k�4�G�����sI�-��>�FJ��0��?X����=�/%X�L�R��0�v
2ѳ8�:�%Z�n'��} ��m�~�}�>I}�\��ө��)�z�>�M�](�<�j�Y���4�Xj3�>}d3��CDI��j,}��I����@��o8�8�dMp%�lQ>�E��hfs��T0	0D�D���K�+��-�m����4���L�>x�e�2n4ё�'�vfG �$\���N7������O��w*�%���j"T��5jj���PlX�H�Cє�� �g��m�IF�C�S�&M�Ԍf�֝�.#
=����<�P^��JE�?��jVZ)Pe����	I�&I@@a�W{t����v�F�����5���'"6�-n���w�m=��En��/B�Ə��]+��V3�a�"ʂ[W0'W�Ц��w-���:��xQt��­g� �-K��{�J���T�:�}�����XZE÷W�h�.���S���7WV_�z�Y
�iyetT��*\bsQ� �-�<����/s�0�-��N#��srI"�( �7Ff�_���U�=�!�U���hp^���4l0B�'<�
�z<'6�(֎�ǼW����k��Ċr���*P&2U��\w��9'
��QB����ʻ-�5BKzӓf@�]��:���M�t
�D��v
�����d~z[��H�6��\ޣu�w����.Ŏ�/��;����	'�]�"i�x�WN+ t�V�>w�4��V�diQF��9�`'h5sD�m~�����E� ��V��&���\oǼ�K��PB���06G[�GC.X��N�d?S�!<!�ͥյ��R�HɌ �����v	��Y�����j�;�"�4s1�*n�Hn�����D�Ŀ�-� ����S+�TFN��$Uz�YѼ@�	���`���)鮳�cb�(�l��hB/�W���Pޓ�F���N3�	@�˿�ܦ�S��O-�JQ>���I�j�P�J8��6ܿC*���{�"�VÎ��@d\r����R�t6��c�D�W�.�v��Z��=��؍4�MO#���@��æU�In��r��ތe�g�<=�#|���V�<��A�[�7܅ t0/Mɪ>���S���ks�2
U��X?(���[���(�p���2dc��6��xB�EY`)J)����!RF�U�|#o EO�x��%eY*:J�W4�H�N�3sj�����%�l�
t5����-�a6�C�7e�)t��o�
C��5cj"a�tbf�@���_�a��V�c}Gg���D��E��B����'4S��U�ݡ��/O��=^{>��8�6K���}�Q�!0o?��53�	�X�o��6����:�rhL5�i8�֋��fRĎ�,�n�ɼ�)$T���q�=۟μ�ν:�K��A���3�,i��н�1�U�Ț�j�o\��~�'V�����:�f����lT���L'���R��EI� �q��a ^Mi��HI��-��%��1��L�+��o)�`7���3�w�g���[B�\s��h����䰣��z��^dr�O�Y��o6wx�dl8ҽ$�ڄ@�0zmr�3<U�O�l���N����K� <��k-&�5Ҷ����Z{�k�{���<ږK�>�Vx��3���/��M*�r������&��r��zL����
(�q�1�Y��^4e�/�	��*��ї���p9���m����z��Y���%u�Ș������Q4�Ϭ{<zJ]Æ�.W��d�s���t& y񽬷��M���B������T����D4A��\Db��Aʊad-��
e);kqJ��]�y�yYb��f�#�I2��ڡU�)��c'���j��H�!0���;^T�0k0c�T�V�X.ǝ�y�St�nf�"(G�|^+kQ�Q���'��k��T�{vN�:�v����KUxe���I����K�����ԏL�ʆ���J���&ŸF6����OS�o�Vnc��4��ք�V^�"���y2��C�m�`E�d��x�C)q`ɓH�DR��r"�&�qJ��献߯cϒ|8�QC0{�b�=�}`K����N����9xG�oK��a����궅�z���b�C��h��p���r�?c꓁⪔�2!.CJ@��NS�is��M��l?מh��#X8��dr�@��m�9�~�V���,n;/�%�E�- #�����4�,�I^��9�_{	�{H�~/�cDgb��R̎:�Ԫ�]TO3,"p|�N��s���̢Mp�h��A,�S�yr�p��.��2a�j�+��>2�+ۍT��ݨ3�ޔ��ŭ.���ܗ]z�$�b������{�
-y���]�i�P	d(�ʻ�[�o�Ń$��	����h+���Z�u-ݐ~ژ�1jVNY;7�č$�ڧ{��ǰ9=��/pz���f����¼�du��kS���߂��x���8����l�;���D2w�쟶��{x�I)�c������,��cJ'�MQ�R�.�kj +�`t��wZ��<}_�ߢ�7� 2�T/aE|t���:�i�~ku�qrcC�-�����}�C�}���fZ%LN׋�)U�o�"��s�v@!��*����^5&Ï�#u"�W�|��hZ���Ob0��_6��Wa6S����o�q��p��#)�k~9^t��R����P��&�\����/d#BtUq�h��Au��S<r���:O��i��4��}��B����%:�Q3h�N�OV�aIqT�Gé��P1�\GbhX���Jc֣�슦�Z�����/�#<<�V�#�����υ�i�{*L�L�Z�_F ���ϸ�����O�������$�Q"3��v�,����|���q�QE�9�~&ی����(�4W�s1m\ᠦ�c� �x��x�:���kh�J�1NK[6BS:����.��XB�r�R�Ī&C��W��,q�1=��m-�-�3I�*��>� ʀ�?&�-�ޑ�#p�$B�VڿL_��Ys����_�?��<Oa�4��F��o���1�W"|~X �W�).Y�g�R�ikPK��`�3Ԭ���xn�C(G/�ң�6p��em�#1?A�W+�0�j֣Di���w�� ˲^f�)���?�Wi�z�C��mU�Ps�\u��_�t�rt�2��D�u��m�_���>�2b{R�B��ki�IeGo܆)��@�$�u+.)���_MdH"f[��:��!��$~l�b�x���Q��}�P@IhT���e�n	6�-V�e�b�?����>1�K�n�kU,���-�:Z+� �J��r����-I�e��^sp���/3ñ�k����x��6 �.�D��u��>s�a?3��h䪿"u����,r\�l�h�I^IF�����[�U#�׷U�@B�:Z E�]�Q�*�{]����*��Y�ź�U�@l���f1��9bᬱ�8LQx*"���/:2�ЬJ��	�)������ɹcqg��؆~��� "��M@���Q2���J�h���p��>��6|��b���[cۙ���@S�"�[�t����c���o{��Q�O�>u;w8��ݨ�κ�2CZ�ӵX�3���(gD��ڽ����uE�����+�����&��B���[�f�cLC�{����zG����J�:�Jd�Dc�-������~�s�X��/@��s�r�G����K�d6�>.��o��q��qb�z��h�	��p�݇ZO�	��}���W��N�5���wn�z�����o�_{��U��V��R�ᯃ,ؖ�8:i��y��B�R�ݠ6��+�{6�nwS��Y��]�ւ�i��ހ�>��4�F�O�9Yuz���v�o�\��suiDðMO� L{N-7'�I$w}c
�X�H�������}z��P�j `��~�L3�1�����I;a�ؤþ^�?��H{ =��_ۈ6[ٕ�1�D�|Q���,�l�J��5@���z��BЃဥ���/�ͳVZ�e�K�tD A�A���sW��MJ��m�� ~��c6�h�ɟ���o:2vV��O�4���T͒"�� a,X�I=��טּ��ǹH_���؊�1��E�^�E۬9�% ����yS_���xR��3|�o_��-�3r)����~m������z����}5v���򺶛t���Dt'l���Ϸ{�e�A��<&5�z�2�G@�C9t`�Y��h��If��o=���7���r�s�k��Z�� ���EcZ'�=8>)�� !�.T\���G�z�@\魲�3�;3�Ȗ�AQˡ���:��%B���@��k؉���"�;��Z��z�ζ�ݺ��/	���J�ol� �/�5�L�K��#�*�C]������cyc���o��#�t�|��w#2�IR��h�	� Ǧ��)�Tj@�VL�X�ܜ�+g�G���,�!]�@�QO�o�U=@5��[���W���Z���tD��P?�/��%f �oNQ\�}��5A�4O[X�oj�.a/'�ے�QG�̣�j����*�?!xY�5S��Cu'u�
��y��Τ��w�X(6je��N��}����ꊗ�8=��-9��~l��ޅm�kn`��Z;�'$�2r��!�<�01,	��+Y�s �ߦ��&�N�!r��Ti��*�F��k��bO~�0��&�B�0B�ѹ�)��~q	 ����l}䌎�ׁF�3�BN�^�"$h>��w�Ϫy�hV���oN�]ҵ
,[ː����|t�W�_[喻��[�r*�uѢm��wTp�ph������}�"gfv�T��^�=Wq�?w�M��5�s��
�z$��ͪ��f4[���3���n-.���k��*@Z�<ec�t)�!L��6wi:���1b۱�S��Q���:��p*�(�2���?�Uɔ;3�����ړV��n�as���N��x�ޭ��	��;�����Uh3�)��LN�}��J���h�U�7`�ِ�Y�����m�����!�L�;Z���U�����;三�2��9I��z�K`���a��_}r:dy@ax��c���W�{OKF2�}r�K00Xp�?T��p��yF�8�!�g�U�Y�[�ң����B(MT&�|�z��[�u����pȴ�PQ��!H�b�%�	\z�rǪ{m�+l��; �fj��w7�%��=�[�;k��.�Mj�����dUU@&�i�"�_��W��zW�C��u�G�w��x1�7Ew��w�=q�'�CA�,]mT���,.�儷!�1M�We�_��Xͥ�C�D� p���L
1���d��t=vC��s,��f��A+�3�UH�t����I�l��~����t���f�b��@P�%ޟ��='��L1�s�^�L9�bh)	~�OW�_�#Mٳ�*��05��rG�R)U���ةi.�\��wD�����!���R�ЪR�(�M|^*���U��+�$#���5�`ʑi���־&u�b��D���M�#n�!�N�����_?B�_�9j�d��Y&�v�L-O��1�@�&�!*\�5�[H�ܴ���:��tN��|ۉ,�:�Y�q���ﯭ͝���� �|�^G���/Ǐ�ด��g��Wǚ�j���-��F%��7��ڈ핲�G��̼�3#JDo�a� cܗ	
8 ���M�7��H˕��ޑLu8���专	[aa����ؤEȫ��4n�z52~���NR@dXE�u��y��]u�d�Vz2x��% 2"M�����&|�h�7�,����R:�2"BX�''���;��i}��X4����Z��5���f��X�I+<���i&�b`��b�C�~~��J֛�{������)�;�H��\�}�Bi��B�Y�c�IB����?u���V�δ�i8CA⋶����������<UZ�@{���S���O+E���~bRq����?�.#�/�m9A�u�ڹPp���H��2�k3��A�?��H'��Gf��|���lmF3�k��_���S^8	G������Ӫ��S�A�Ω�Mr�Yȗ`�\<D W\��d������-\	�$�X�]f
z�u%=�=�0ђ6����|P���|�9qypvU*���q�여xx�fs� R{�^�$Σq�f�P��#�ݐ`�X>8r����Â���s.Y�Am�YC�X��$�"�$I��a<9�$N�^�ZG��;�	Y�w����ޠ���$M����i~c��RQv5;0��s"��'�T���.����D<^���Bߣ�U|~
��?���[͂dk�!��*�4եLyG�%M�|/���#lm�aQ�p�;��'�@�SY���E�D���.���sǍF��U��j����1L�+O[��۷�P51I�lL�����1��svȰs�d�lh$>�,M��0���;�,�Lz0�,͐�th��'г8&ˢ�B��YL��g��jsm�{��4`�0Gd��> +:�ł�sDZ 'fۖy�$�Z���s�M��=qO~����j �>k��jq��X$�?�?2q+*��ė-��P�|f� ��]��}a�����#�)��q�� ����`�r���ot^����k�G�w?3�ToV�0d��0��mG�~�P�U���Z|�V�k*��uB�m�/����48�-��"6d����t
�{�>D.�hfOv��4��$��*4��m���1��r�|��/���&e���(&?X��H�!a�݃��Y��i�k6DAO���B�[����ǚ�`)/���W�M�|h��grS9d��_;ek�EaB訉�P��}�K�Fs��3�ʩl0Q�9�*�Q}[�n�{�Rj��t*9&�C�%�?��S�W�3�?f/�0[�zq3�@T恵f����� �7�A�u��w6ܮkO�@?dK���^�X�U&t��"cB6��՞%��	�D����������
C���,e�M}����/�T�ۅ�B^����Q�9�v�P�Y{ܱ2�e��4�:����T�>scA��93Oڲ��Zc����>�^f?����0����w����I�a��7�͉|W��\`f�c�ʎ
�����p���J!���f�]e���q��}�G�P����)��=C�!7�=ki3�h�r�#[ ��5Р��=n8ǈJ���~-c��
���i��ƻ&�^��ӱ[�Q��Z�T5�BhI��^�ܱ�\Z�쮾�0�%�"%ȎJ_��bY�3v3MP����B��1_�y �E��{j���ݲL\Fd�p@Z��>�"����S%6�R!��ns�3��/�\���O�hiL��Ǹ�Ւ@a�Ȅj d������e��c'8�Y�T��"A���`®h�ӆ�!�t�"���_�?b*_]���̢��:�V���N:�Y�v�"Q�/���lc,��W�5�$����0�[.,GbT���a��u��KLx.�'S���M�� ��{�{O��=2�a�N���sX�~�}����Ą��fDT�YYn���Zw������tB4��4�nh�"W���U���H>��j���˱���9rEk���P�-ȼVz��ɉ���͏u�Xe�P/Æw��j���-[b8E�c 7ޕ4��3�z�r}o�P!�0�١�MY$�k;�����S��� ����*pݗ�{��T�Yszݟ˛��G������TG�;�8 �JQE�D��/��r ����ɉ:J�e}���g����jS�zH}؝u��V*���Ar��}�ً��!���!&\A�����2���K&��a�Q|7+�β�]���^_9�<)���ʥvD\���r�Wv�>�g�q�/`�7��\��D�(��q��`N�/�uQ�#��_�9^�XRЋ��7�^��2Wl!Ӗ���zڽ'v�-����A3����[�������}h��]�`�N�O����pϹ��[��n�@Ws���\'�X�N��};�]�m����q���$�Go�3p���j�wO���թ�t�m�}������x�%��R8�%���)�$wA�/��+y�����B�h:E,T�]��<\�*W��]�M����e�j.�yx�R�h ��+�_w����`k���,HA�����"���h����@h�&��ɴ�Y�V}6�KA��P��j�[�J�&5��t�������S�:�#Q^���P>�`���X`�!f�>0Țˀ���M��W��2�)���	5ָ&tBZ�!��p�3���0�e<g@,���T�'�GA��t�3�9�74�j�����s߷�m} �_߄���k�qq%͉��K�R]�*�-"����5EٛD�M�����6�6]�WC����������$�1���� ���cx#�h����҂��Nl�e��(��X����?���|�,��3�ڋA�Qĉ���M8fׂ�$����
*�Yz��S��88��*z?G�$�V��5��hT׀\�B0�W,R�4<��R��&b�G���"5�'IԔ,4���_�D��(�,ǊUlv�.G�+Mk��h���Hܦ?�#B���±��d����W<��w�v�Ӏ�����*�ө��tv �A��Yu�T�E�i3��Ȟ����G[b$M�o}�]+Et�=c`"u�eo>b�n E
`������L��i�p�D�b�M�O�3x������p"Ȃ����;pp�i<4LQ�/�o��@pq���1 x)!qN��`�,-���Yf�o5��7H���@��̀�D���Ȃ}4�8[��֡-��v�z�n!��Z�m��\�.�0]���>k�b7��:dR�l|�CV,�� gv�����&M�P����>��p��M�~�[(��}�!磽���ʓ������}�:���a��N��܆�K�d���A�� H�I�ڭC�7B9����'>�ɨ���"��+t4�SQ�ź�
�[��W5��� �ؔZ˱6鍲�c��9@|M>GH��w�C7y		LoxDT��.��.@��O�b�����=�qN�z䂟���믿ᅃo��y9ȗ�CtNH�n ؋cIjZ�]7��^�;/�����0�VR	˦=k�<�tF��z:�{Ҥ8 m��-���)y+�Ɇ��R�D�D�A�Fyq�����Z������!���'�@8#7/5iI��As���܌4:����t���R+4�A�
xğw]HQê��3Ng��Aؙ��C�r%!���pX�y�e}$�Ԍ�޼6�F�ǜ݊�5��o���NU��ɟK�0����̠��C��:3��Ζ%Y$8,̺��Wb��T��{?��}|��c�sq���Hzb׌��{�t���1��%q�_3s���IN���ÿOp�߈/s��O��񎢊eLKg��8%HX�*�J��wd���R�k�S��:(���j�i�=��h�v�u�����q���&�
��Jj�9�Ke����B��ڳ����v�Z��ʅRg��	�9��ҵ���P�]X��	��+�2@����N��D��C�Ԑ�.�z��;E��]�EJ����B*T"/�&hj��my�c��ו-��<�'uTcģ>��,�aw���vh�����j�ru}�ܶ��9C�h��?��,N6�t���t/Lz�"�!@&�v�'������M雏k3��/5O2���O�G��>m[N�g�DZ`$�-ӥ��L6�h�;&��=���7x�Oӗ�nDj��f_%K��zy���TB�sA ��+�9���$AL\��������������#~D�bA��X��,Ok�?t�OV�q��̀�׉��O�r/�9,Ս��+h�M]W:����.w���[�<�6������Q4x��>�Q�
cp�Y�Y8w�o2Cè/�q�D5�^���<��+�2x�i�#?��3�Lz��F}oۯ��T
?����%�=�'�9�p����)59����Ù �.`���SP.H���+�c��$-�d��ڼ�s��H3�'@Oب��U��+�t%A�C��S�sr����$y1�v4�f�XWj����,*�w�F���]���F*�ͷ~&���D����	E�t�)�įMfQ�H��.u��} �Ȁ�����������ҁ� �����.b.���X�,�u#�|�N�{�� T��J�O�����ϖ��/�G�$�I���B��*e�X��Xɟ�D��W9�U���:y �vŶٴ஠sK�:�7C��M�4��o��QҒ� ��k��v>Ӗ��l��������"標��}�&�Z��q���'�}%6k5�q�H�O�DO/�I�N�?Ѯ*�NzDE���a�h�����6Z�*%�� �0;|JIX�������/c�Fk��m���?R03gK��� )�)H�j\9Q��Kȏ=�ƭ߫~j|ol�ךVja"l��6��ݪ9g%Ij�Ԉ�,�!�ቢ�J�B�yj"�Ҧ�-�pm+�I0Q�fO"n�t�To^?n�Э�T�<E�je���S 0�q]a�#@�G{���&J&����+=Tz/#�������D�l�"�v6�ϑ�Ӭ���&o��\�Pn�v��~�Ӕ�@���b�h�b�詀��t
G ��T�����ݧ�o}��9h�u@��m��Ȇ�(W`b�!�z���HUv�غY��CP�%��7Ҵ7Fe�e D���)��izQ/vf��@�D���QMVQlbБ�W6>�5�l�}?7����	����6\NcÜ�Vf,1ȸVRbJ�p��Yi'C�E��Տn�8A����8J�n ��X��	�a&���j����������J�[�:�c�:�����D�=��]����}I����ޙ(�w�Zt�f��4����ܖ$S�@P馛��f��W��'��+�����<���=�g*���en�V�����;m��6�.R���U�����x�����1t$����ڱ����2),�f�t�6�2x,�9�V(ɹ^Ѱ-�����OU�ߒ�x^�7���uڔ��(��� "`Ӧ����c8�(�@.1�Frm����"�,�O�{�8}��|FJh�iӟ�J���G�Z����Щ?��{Դ[��M�Ҡ��Y�S"F
��\�A�4�I�8˰<�C$䴲�+&�}��('��\�|\20�%�[�}c�q�?d8����v�c�(�,���	MR�φ�$��7`09}���,�]褟�dI�_��e*��R՘R�1Mt�w�O{{�]��4��SVυ��L��t _p�=��s�*]��eGx����^�h�ޑKM��}���1"�09_0�8ٱ�2)Ԩ�0�w���W�A�������L��������O߉�׍ɑ����	!��/�Y�޺gH��fmM�[g��2��W�ϗ�2�SG�'��_th~�h`�L�*mɶ�g	<����i����j���s ��	�� ?rn���㍁QT5KeZ�i��8n��;z��p�jp��e2R?���H��.�,��D0*97jzm��QR�ˁB� � I�ۄ�6h<����/�}>���F�뇄�M�\�

�6�2��,�%%'mBC���؈U/}2�Z�]M~>��myg隡��E��gD��*pw61�?�ú���u�1izq���ꦬj�8!���8>��*F���?�7\�b�PQ�.��?�AY�~�o���`Z�j�Z|J���k� ��$<y�2RS'J��a�U�'��+CzAȺP3��t��I	����$;��tf���	}M�a��YO�W��+�su�r����:�����}po3�%�BPj��`�L��3���`.&�t�y�Sz��,���F�L`0@���!\�0��.�1�='�{�	��73q�/�Q�]mNr,�4֯�qw���}�=B}|��4��9��KV��OD���.����[sSb tVq�{A�;n�S>qL+��Ʃ���BF%&4��`,����{�ٗ�U2s����|Ғ3���0��}`���x_p4��E�f�;��Vk$�b-��e�f��$����BG>%���,�soP�>E<��f�hkk��m��%]9����C��*��"�?�h��b d$�u�Ӣ[c)�S�ά�_I���i`�5�� ����"��V[�)����ң�f9��3CR�g�^N�u^N��Y>��\Jd��^c<�$w��咞�[�`ٝrI�2}G�jAj;�P���U1���=�GSK6ʃ��n<x��'���ZsUf�rvU��ob3!v�C���k�\F�31zE��,�F�ʾ�zp�-�)J4���"[��gޑ��zr~`s���k	� L�_h�C�~��aG8�a����1���0zn�4��S�IF��!����o�6��h��y}�%gv��X
^	�G��ORZ	��jg��pq���>NQ8T�d^�Ahn2�q������O�1Ӛ:Ȅ�uO��<4�bi��i��+6_���An4��h�������/Ñr�(���{F5�S�x('x��:@���>�Z$Z�s:T��.����f�2ʢ�)�ߧ��2�JJ�s��-2]ɇ�x"��=��l�z�5Ya�S��uhe����i~�:
�F$����S�V'��0�|;b�C��(ps��G֌%-�.r��|2���Mi��Z[���F�QE���ڍ��)#*�u��Q��Y緭~���!u�������lnJL�)���G*�-d�ĈM�5��s/"B����?vi$|CD����:Z�!=���f� [�����/�
��m;}�fw,J�'��60�3Ѓ,';�8�Ck�LHLi�qw���g=�W9�x�,��c���aރ7
{�hYXI���d�*ٻ��-/wܟ#Fb�I�Y:#s��M�����<������������f��ZM���GJ�B�l+/�!|]�q٫�*���D�.ð�FW��zj�׽�~ã%Dڸ`ӷ�]���@Ԉ/m��[�&E��U�v�G��\�!4��W<������oadnFA�_
	I�R^_%ar���vv�M�~H�1�[�ٶ�m#��e4Vy�,�Κ'���!�d��Q~T�֎
��J�D�h��r ��d�N�ъ��]�p
+��VU�i|��|�w{ ����&�	>�]t8��c���6b|;Y�"��
6sk]iߕD6"��z�]d6Yj�rgZTJK��Nm;�����Q��K�����af'W��R���&PE����=�Xb���L+V��s��չ,���"<�CAm#�vEQ  ���~V�\���Y�����#����{�&l^
�`>�� @BTp��|2���FO<[ˣD�w��{�e�p�^v�)$
/�0m[2�~�k���p�K�D]�R]�����&/�h4Y/���z���Ε��p�v��t��>����Ő`kTk�z�!_�~l��-����D�g�{�C&����Ǚ�p�`�YF���v~�H](�hV�A�Ϊ�x����q��S������C���)'��7E�,�^�&��0o��G�+^�)���~�Z���<�	��#�H��p��f�Bu�#�!s�X��=�!s�g!U��iZ�'�e0�Q�����b|5F�^�mX(�TI��dT�o gKi<������_1l�p.R�WU�!o�v�C@���@���c$81s])��S�6���$�����BZ
�<y�uE+�s�B
��b�O�y�ׂ�55���q,
f��za�P`>>u9�|�N��W����H4l�4�:��}?�B7�+�CY���������e��r��7)܀�?_�p}����peP�9�k\�'�t��M�{�3�������b��%"����/���H_��u�]��g>�f�B1�p>?߭�4���p�^�]�H��f���O�°W?ͣ���T������]U�P:^2@+��<E�=	|u3B��	�g5��j�������XZ&�o �=cp�/��)�1F7�Ab�/��t�#l^�`2�1��{������>�$��U����^���z�}�ښgE�P=���Qr5�ZV`2`�H쨩=�/L�CpkK�*����-�������a'Kz�{6�:�#up{5��;=DfH_9M����4�E���Id8�o>5�>{�{���
+5�=�����e봋5b7�C^��h�auӋ�1�n�Z�tV�`�A�_,��u��K��^2�'�3�֗L0�H��#�o����k��@}�X�����Ԍ-�g�g��v�ã=��y�l�>�A_��1��A+��D����;c70�F'{p���7�Ze������ 16
�aL�f yn����ׄ.r�S��FB�"ڳ-�BW�ή�a�xN�]*�ɨj�A`?��ֈ�����ȷ���}��LM5�����Ѝ��8<��9Qܸ�/�-��HO#��9������ S3�V���R��ҳhhAb��|-<y?ȅ6.a5;�3Җ�:��7h0W����X�rb��n�ՠe������W`��P���F5q���r����\�Wbh�$�K���C�VhĹ��>A���*�.hU���X��޽��d�><w��:d
�Nɭk�@���Çׁ'����Y�p�Yh��Ih�Ҩ�>�;��^�¯��
���{�>�m����]=�*<ԡ��~b�J�����$�n�yz�k�o��Rz�bz����O�~�a۶/�f�沗���;�9�5�'NO�֢N�K��KQ.��[F�މѥ��/��H�vY�I.W=��˪�k��8� �X��N4tI��k���U�͖fu+?A�K"sg�R��܆H�aД���pLn�lJnj�jYG"���(�t����,ѭ_"�iK��q����6Z���H�ɷM�R�L���H3~����w���P
^A��z7�]!?�3���d���D%Tߢ�I�̠c�-��T�	����ӳ7�ӛt}�]��_��ۖ����_7of�_Q�Y�`�q!�<��
�2�4/���%�jb�q�9��%���/�+faA :!u�M��.��*b���;ܥ~VU�z������?OA�RM#� %B��E����9�Wԛ^��~����UG���s��"a���x�ZM��P�
�Qظ!��={����F���Զ����pC2������S�����#lAS��I�G v�',��h�+�~G���D�a�BF �L��%څ�6;�	?A�f���ȳI�!(zG����E�:3	2���R~�r4�޲���T�H�c!x��".5��e|�@��Ɍ���I�m�<�t����A�$9�z���md��r�eaT�?_�*��� �~�^�Ƽ���e��_����-��t�w�X���?��`��u��l���**���
���Z|j�Z`��{���{���r��'�b�Ƕ�Y�d�ěLd?t��|�>����:8��K�̱YUW��:U�#�T#�A�<�_�@ZY�4-ɫQ���цf�{(�� r����L�d�\eN�T�e僗��{b������7�k�aӶ�9������C!}6롭�θ�X����t�Y"=�����>�' ��$�/|�n����@Vf�=\.g3{n�z���Ə���2�U%/}�Bؖ�S�eY�Y�����}��[x./g�(mZyz�@�/,���?
�>/�.A����FWZB�hg埠K)��E̦�x�EBV�����-�-r�E�o=&���#NR��H�u�W"�b�T������0 �$������+^/~?�a���4ʴ˞p]{z~���� ���#�J�Z�e� �>�Y�ݼj�8�Օ��x�)�]K�EP��Rdٻk��,Ѡ\���n�ЀP�@`�r2Is I�R�,?g�[�ʛ�]�h��#`-'+�U����üQ\J�4:BU��LE�9�o4�M�{N��&q�D�TJ�&��E�PX#���Ç^3�+�fѸ��?�	1��U	/%l��?��{�<��BU�AŖ@E� ��#2dK�R���$g������1��+e��|�"��R����~�烮X�`�h;CĶ�0�*ꅆ�u�f�F�0����V�X� ���z]���W�pFNwD0���A��Ua�u�d��ډ�W`�wG�V�S1P����î�J�J��B�����g����8��߇�޹Y�X��nލ�bͶ�[�g6j��J�m�sb)D.��s�5V�*xF�J0$��e�⟩�p�u��&Du�4М�!=�<�)�g��`M���$=C��A��iNW
˿�8��ŵ�d���Rd�����5�.�L3� ٭�|��@PX�*G�}��9�!;�7yG��3l1S����L,�� �5���'	��:jk�6���3���K�R#��v4V��e��$��:��������$�-[x��Ґ �z�*�u��}���)����Z�qK�o�dO���ӓ��,�W�#���3��)����P(AxK���#L�|�*���N_�Q�L��yUƻz�oEB���~�:r8@)�8�&���Cj0�.�A�տ�N-6S���1������|�ah�C��1�e�>�{X���;e�7�;b.{��A�`kZ�lؓVC�s�6 xѯ'qZ�x��u��(�*��Gvݽ� �о���m2?��ϗ�W�J�hAS;v�y^pͅW	+ҔD�b���	�z���^֔��G���2��g���	����^<3O�@��{�y*�Rؠ���k��3Q�@�+j�G5q*~����y&����\����)��%���*��Ez�,�#]�edKH�2bflD�r���ޟ+Z������!i�$�6)��|-]�=}n[R��\h�+�p�fPq���0���yQ�G��zX�`�5o�Mb�(e�F���`	.s���*�rrQh^6���r�|��HI[�q ��F���%�1)�2����;��0}���쾹U������n-j�j��9������x����_�~Ӈ�R@u�%�!K�r��0��qۡ�X���i)d��q����>S�L�����)IZc}n⣺F5S/�����	�lVt�h��iC�2ox������ϊ��%� R��d\�h��� ��)S�4"0��՚t\Zm�#������<�nc0����]L��J���w����Qz↕�b6]�ں�ɪ�q� ���-�&��g5з�p,�Iu+���2�PC^�Ń�����10�ڹ����]�y ����*���=�tt��C�`�vJ��b��A p�O�rX����	�{|YlѺ9���л8ךhkţc�G��f�8|�
���zW'F���b���s���I�Rz�)�C9 TGo	m�� 7�����	i�L� es YYf�<����Ve�'@��L���">+|��+���k�q��ٓ������c�ag@O�ԡXo��r���B�;�����aw &
Z~� �X&��*MB1��G19Ly�2�[1�f)whnC,��<[��w>d׸�5��|t`��z؂K�L��ې�ѧ2�� W���b�Q��eϦ~`N��D|���E�'���s����e+%��,$��y䒨7���-�*+��c�C�i�6����/{�#ׅA:%x��/��]bִ�i%*�u��{�Օ���0�1��kJ����t����5�l9�r2:�=B�a� �Y���N%=�p�K�Fc�*����n/}QXN[hjV-�D�x�)��w�w��P����M����dF+�U�
lf;(s��&�Dnˁ�7��&D�w���Ѝ�˝D�J���w����o�������\�G��`'xZ�������)��C��)[��JA{ݤ�'4碞�N�I���8 ^�v5��-|�t#�fCAd
Li?}-9\x+&+�h�g-�=�}z~��q�%�nՐt���f��@���W����j��-�{�)�%Ɍ�Ā���J`���-�S�Y��ư7�Al&X:�kp|�X)���J��k�w�U��r���X����Z
��o�¯a�&kB�&�5�WO�S�K�dCV�N�Ƹ�1���蘛�8J��H~�JR��|��_H�;�������U(��'H�|���]xp��$� �8�� _E�� 8 
����O���Q�o1�i�-�Q5n���ò�!�`��d�i��W�#��U/O��(�1א'��*$C���)�A勧�Պ����/��ɦyTs V�H+J�uG'a���ū?OSe+�U���A�c��5�g$ɏT��T�w�?L��CH�MKź���v��J��A�>+43cA���I1��=����..��;��@�~�l#~\I��{&ÃaE;E��t�;��>�%mb��G���6����1��uD�,�鸔p<m �F����5XT�tl�z���B~�<�~3zˤ�o�SL�x�:,i࣐�n��<=�h�Gf���4�j���~�8w�0h��U�L�;fr��D�wع�/��C�^g�]��q@���+�NX#��3�@hr��w�vi�?7�P���o+ش	Ͼ�ΨE�W�w�t�����[.a���O�lINH��W��^@�y,�j|�F�c=��k_Ū���a�Q�����C��6>�ec=C��'�{�tqL��uQgd�*%�Үa��iOf4rG�z����*��Q���Ānu�ab.�4�Z�?��_���Ɔ/�z&����}@��r�:W@Xv�߄܄�r�n6c72!(�B�+p�6v���3r�"����n+k��T7=�u�/u��X��,����m�1��ff@G6�R���{�?��J쮕�O>�M��~nዽ�l� ��q�� ��c�l���h��ݢ~%ź�I0i�[yr�B��>���[�˽�^�p���es=�>x�v���
@�l��Ŵ��as�#��'y�*�I��o�8.z˼�"r|.:�u�1Ӌ�~'��&�>�t}}��Ԫ��pW?��,W��[G�����p;?R�ꅝ���K0�}�����}�����O��xR��`������VP@���V�|����>�o�sx�Ac�3d}?5�D��Ѻ��N� ��X��y���*I�g�n�)Toy�wV�M�)��]��5��GXV#�Q���Ƌu���6��]�q��1���S!a|�^�?�����Y��6dI���/ZY;Y4�l$�tv�5E2�������Z���A�/�)e���Of�v>����8DX\F�N��Bj�@p����X|&�7�?�b�$Ld;:�/j�D 1j8��$bC2�<��}fC��KP	;z��> �혽oB�86x���v����u�=�Ū39盗�g���(�^�@R�ѳZM�2 )�b���t�+��#�,r�2|��޾H�i�B&�ȼnTRD�/�F�"���FpM\��W�86��m�Hc�"W�f�{�:���M������T��U��z����ڞwVZJ&�Ω�L�(8@���`��a2x��}6�m�yڷ�Њ��a,�;C�q�y�X�ъ
u�g@������W9 �Y0�<��zH0uR%�C��z�oC�8��)��,G0���6�>������E�ɧ��10���P�����Ǉ��	]"Xp`7���|r�bdM�Z�{WV-qx�Mm�Qh��RY�ahm��o�	�ٮ� ��Y�v�'`e��X��1ꎰ���x�h�XA�"=�?�Ópђ�Zò�~^/Q���:�41Ii��Kk!���}���~�W��`E���[�:?�\��,���4�55�휣	:۽$����I�qKuW��1̟��8ᒈ�ȕ �o!{�$����ҿ.#���­��f	N�0%⨁3(8:T�\�^ˡ?�Ew'V�
b#��C7�!bz9��P���$�D�4z�}Ԫ�@I������F�z�rE�G�����ی}A��z����\Rh��z�0>�h�z����cYLI_��(��;�/aa�.[CM�M��=��*dB�E�1�%̴���?E������z;yJף{�<�r����ϥ�;9����[+_aY]�~)�C��F�y1�X����X˗��.�hgg`��a�������\��qi���������,�D�0\u���.����&c���-|jly���o-�~j���C����;*����}�ߤx�Fe�6'A�F��<��"��WEX��}5�Xw��	||�����##g<,���u��>�=��ޕ4�+u�^X�mEύ�.뒄�Q�v/~�q�m��'�Ge�^�0�@a���l��e"d9J#��z��㤅0��O��o|g�,����UotF��;�Z"�k�%3��%��&&�����w|Л9����맭�w9oi�ؿ?���ݒ�]�b[�ᨷ�Y��4�6�C}\�_��F��ͧ�|����)��3������Yi��N8~횞_������3�.A����e/�/��Q���
I��T�X� �$'�2p�J�w�ɕk3�IQOܮ`�����[ȓ���ݱ�M� d^w�l�g8�\� �LX�f���h?���Nh�¼��w�#�JV.��É�R�&T�Zҽo�js� RA�'�����wR�����;E����ߛB�S>]P�V�{:IH_�[K|d�J���vB�>G��=g���p�Y�3�͹q��P�oO>g�rLT�!ђ�o��ȣ<�G�O�(zv���c4�ᇮ�ye�	����j1��)�f�����Ũ����5»&�A�I�9�,�Y�]�	B,�m�O]��d�^�櫓�%A�Rvıw���;5��ؒ�^48�))�*����^���/��O��	�gm,U��F�=L�S���q�I�6��V.%���PK�&u8rv�H͒�Xx�5Q��2v��J���K˩D_t}��9	��kv��X��c�C.u�W�+����� �O&��X�c$HBP󶱹w�2�F��S���o���龋���G�!���e��35�����5�hn�b� �\�/6��p/7��?�Ph��;asrI=�,mS5�(�Є�h�V(x��8dʐ�<��Ys������r'<�����_�g�M�?q�O���{Z�W����7����4�IШvu�d2�	�F������Z��a���(o�7����DJ��V<�^C�Y���|�f]��|\<��2Bu�x��<��0h~�Z,��=�����|�.����������h�m�Ei�E����C|L�-&nvV_ԾoUOw�O�B��J��l�7�I¾�oez�-�4�U��q���rk��D�S=9Ւ�7\?�i��y�?�v��?��;�G��rMtLP^Kv�zp��&<������(�⅘��*ϡ��:�#��Q�;�QzS���>��ǌKUO�԰{�������q�����73�hW�n�+��ִceb��Q�&i��6��=KIi��p��)��	%p1�%Ͻ�����+�g�` d�?�&(����G�-�ɱe����Bv�=�Jc������З�fZl��b�ص�� Y��A����ʍ:�B�*}<y������X9/M��Zج�e	�So��C%S����+��
X{�ռ5R���sf�P��$VS��X9�PUۚ���7I�I��a����Һ�$��\�ǒ���>
�)45_q��Vӗ!M{��	���7d��w}�=��p�x����|�-S<�����٬^_������eL��x����+_��N��hoWV�'��4 ���C1����!t�"�mV8A���hD�׺a�$A�wQ�U��Ka��[_����,�C���>e&'i��ٰ/Hf/��C��q[٭<�q��=Ձ9q��6����2vK[��r0p��h7�'[!�Q`�h�퀳1ZJRQ�Fe�'��f
g.|���&Ф&��.wߚ?��4 �X!�*�Q��G^B9n��3���z���` ��A%�,/s�k�� ��%�Eq:1.I\␛�A���MeQ���iZ{�E���
��~Pd��j ~�<�T��?�?-\?
}
)>2",�k�.0�+�����ؓ���J�)��=��H�wF �=�{��4�P�A=n�		R���.�(Z��ޥ�(���7	�a�E�+b�`-V��V��w�������=�A�z��m��1�b��� �O�d�Tn�b�&��D�J%�#�Dcb��T�J>��z������C� o�v������9�z���xo�᷹��F}�۫)��}���P����H�����#	�,־U5�6!R��Z�S{��x~2o��<��d��n�+8֛F_�u�.m�NEz|e9fw��<���1$@?p���֝Ů�1�@`��O�L�ԟҲ� ��� 0���U�Y���2��a�ڞqv Aّxb�d7n�΄�$�>�q���s@>TEm�i�R��g�"�-��sF�YnX6z�wB��k;['�N�_b2�%�h��K-����;ǋw��z1�3���FKcp�jɴ}��3!=��F%v���c��?k�\�WdS�"�����2�b�w��V�O�L�Y2)�p��`��ĳ�=6E�Ul)@����$����P�>Y�b���(RA*Kx)K���[f�����T���pX$N}�c�lf� �&8��EJ�SP�m�����~f�8��v}n�,)�Eo��w�@�sH����^iy�.�ɦ=�[��^� *��һ�:M�VF��V���Q�-0J�s��$��9S�w�)b��W�ćۆ���}�����J��h{�)��x�����Z�.אf�R����\�'�T����<��i�~�DI�
�w��;T4A���F�>un~Y.��쏭���U�\��}�(��~�j�C��;ڴS�-�c���4=���s��?J	i�+���8�Ÿ������F��;�������9�����	�͐�#7F*t"�bDP��+��Ho0Z�eY���<昝$ؠtӈ�輸>������{�%����S��=�q�C,"�毇JM�)�<H���~^�}o̠ͪGp��j�28E�L��s��o&��Ƞ����`0qR���Qu�{�$�X��/9��E��<�.��0�Ԗ��Ϛ�H�\��L7ab�_ /߽���
ʏ�OK�
0�i{+�gU0?QX�$�o�q`���h�F1��w���k��A�c�kۋy����q;�hvT��t��E�V�g��vB������T �!�LZ�oǃ���㺿��>�J;�K�b��1����b���zFM�ታ�_��{n t����*M*F$� V_}6N�9��L���i�w�H�:��TǇu��%���+��E7U�t��'td��+�td�ӯ�ڷR3�x�;���w ��0Vm�M���;�?�Sܢ������ePA�wZ��'f�d ��][��<$��Q��lq��Ш�ɪ4�x��̿"y�7�ww�8���$�n�¹�������XG��,���D�A��`�G��YY�X����b̴_F&�M���_Z�̻c�җ��#�lUA.�7���c�so���0���w �$a|KK�'J�8�$�j��C�����fkƃ�l���d�5$����-�-/\v�	��5��P ���Lx)��*����g]����wΕ��5�h������+	��pHM�c-���F�	��{�<�Dy�k�$��s4�5�2�,��W�TR��E��L�W�~1��oW�5�R����l�3c�M�VM9�����4�9"՜4b�h�z�7�2KV�]�s��s]d#���F�/��>�����Sq���[ޣ|�T��=|���ʲ_��1���nS�D��sTX�N	b�q$i�t#���5@k�{�I�Q�R��5��"V�|���:��JQ�.#��{og�&�X�,8_l�'���@!8�)�\,�7E��!����h�ע�Ŧ!Eٙ���mG����I��llf����j�_j~�TX�3���#�G��?�NJ<9Ň�os,�/�ԇ���6�T�T�/p��K܊�M�!1u6m Y�r�q ?n0���������X8p4�"��a)d��De\���}"C��4`�S�B�[��.��l+�y%�C���Z?h�t�.&RϺ{�Bi$d�p&Q������t��г,>S�N"2:���C
�/Z�@�e�R�q��dJ#'�7���F�i'���G��u�	V46ش��#T��qY�E���0̜�r����٣�d���{e����N��$[��У:#�� �ޡ�c��~�:���l��!�X�ͮ�QZs�:��}�3�9�i_�*��:���
c�9~X�k�ِv�b!E �����vQ��y�+l�P-
�|���u���v$/7�����������o;u؃J{�V���辅y��dbEa�ss^��E��&��h��t�͍+]&��;��y"N��1!M�`�=���v��%�#����Q�	.X�n��v8�1h��&r�y.����E�����LX�tߙ>��#������W ��A
����_�N�R�	�?�E*J�,Hl�0�-ű@�׭��X�q���a�W�*���>YC�7����Poi��mژp��ìa����G����I��ͧ6m�B͞�%�M�ߐ�M����b����-х�1wӈ�Qi�H'�h��i"�����o��K�&7�|k��b���� )�mj��-�ژ��vy�ʳ�[)�H��jǧ��+�#�}��J�����h�'�{������}�.-��2n�fs��ɭ����K�4^^p�*o����nm��'�?YD:��>ѱ=��2b�a����!t{����	�]hԅP��:�x�6G�8��Q�>,�W��Qt�)xQy��ꋈo�)��7ѝ��|�\Z�0m��(�Qbj-��F��>�pUgt�ķ�O����@�9h[�J��]C�Pu�y���;3�3�bW�,#��kM��[�0e}�Ao�[�B<�]�_�GC�hl���o>�ǀq�'�Bl�ҏ��^�2	Au�yN7�^B%x 0��v��.�|��1|w������L��H8�K�t|�V��Д�(��dS�|���Ѵ��y)@���=h�!�-)0�iHv⨢C,2T�2;����������U+��E����jHv��
Q�;XX�Kn4Q��%�Z�#�K�3�[�ۮ�BֻP�V�E�����m�/���iL�8?��8c����������P��:�M=��p"|l�"쵵4��6݊�u�1�k~�$�	?(y�v � .����7.�1�ܤ-�DRZ���#:��˗��M������&��B8�e|`�b���.	i!�a� a�`]��T��ڶq�7��"�ՌL Y��IVyC���w+Q�;U_�V�YzgT�}1Bz��5��|dFҩm6��
1�1;:ű+C&`����d�1�,�6�"m�[@0.�x����IsyZ����d �B�ͩL7 ����j�%J���ɻ`��5���"�Ux���g�Ƅn��b`��R��m�x�SPl���[�%6��XAC"��h�ǆu=�t͢u�&��w��i�J2���Ά����#KWi�Lߎ�G	��������t�pp%��6����]Z���Z�ȋ��~ �}�W�z�zx��k�e�V���a:.�ǃ��9�]Pw<=F_h�C��Aovj�e��	��R.Z�A����@�a�(9�[.�l�>�"�_��=L�H�h�������Z�Co
L�� U���Dhx_U��t���W��Т�M����+�ǃ�L�R>a�ږʝ�
pB�8��kԿ���v����ַ��R6?�^T���6��_�s�Qm[�\+�m+ swh����v�T���=Gɘϐ�'��*!��st_m�2��#(o�;'���D�ߒ����Gu�4�U3g����z���t��rn%Dz.e3�]մw���L32�h�����ܰ��i��5A�C##�e�T����i���r�W���Y��
m��^���$����~)��;^�"�wi�/<ǱU���7�����F{�h�A��0�mA��{1��S�����b��3��sZdf��L ~���ht(��"T��WI����^�m����r�&���Y�5��b��X%���`ď���k.�OR�|�Sx��Y7��w����F�Mj�!re������=�Lt���A�r���ɘ����zr5��m"��c!�Bw2|ȡK�=��Z_�i���ط��]��ǩn�e�	��)�N樫�Jh�4��B��ZK�Y�7��*�((�� uدm�1OQ�<wmq�i>`��#X-��z�q�v�)ui�b��2�1Dg�N�'���y�9�Iw�E���Ğ���.��{����͝��ʤU<ǔy��s����K�V�
90��NC�琜�b;��[�شp�|3i0���V7����X��_�e�J���9��f��n��I�J_1�J�wԂ�$�\y�0�h������Z ��~e��<@4��|)3�.,�]�L�=zY<��Q��t22��iR��T���gߓڣW�U�1(B�,�M��*�D�����>�G$���{`�(�m~���s3���0���.0�q>��j�uߞ�޼�wy�S٠��3,Iv�+Ծt�d�y@q$�8zKr�J�m�T-���HF0v�G)<)b��� _}�n`��XT��L�-?�G����{���4��|��N�"�R�e��.�=�"�,�2��{�A��&�-�r�����dU������7���(�5���Y��WI���z��8~����e�c[#����/Aj>m8���U��7�1s���������V�5:�vHן� �L� uq�6��om�z�"Fߐ�Eu�,�[ z��B���������m���/~�k�`�����Zͼq�63�������Y'�&vf�Y
%�w�����#0H�ql�� ǧ�����0N�E�@��̗�=8�K�U�4p�ZrE�fI���y��P�Q���T���({n�ȭf�&5�J6��i�������_�x]�5�6�1�K�+�?C����&���>y~ߦ�Eb	I�g4�NT.j��T��"�ɐ��a���Â�]�Φ�02�����vx=b�37w2�]g�Td����n�f���mZd��b�
���8I�y�~PH�	��[b�X}4�M%G9츅}7���/at��A|^fw�h92�����w�<���b@A�2,h��PfS�;���wfx��k� .��XO��H�q�������PZVW�s��qQ�i1)��I�Y���f;��5��@�Zo�t�B���`@�v5��N��1J��Fzm=
��̘!d� =�#J��$b<�V���I����f9?�l%@]o%��1�����IhnuN�Q�a�lhŴ�_F,o���l
N�2�"5�y�3��إ����Ȣ��W�#�y@��[/(�|�����Vӝ�!�C��ƽu��J�p��TL	O�"����l�v���#w��'�#q��A � ��Iۍw�,�~2�>0������my2��VR��V_�-���qCaІ�/�`�
��Њ��Je����1�-g�$�,~IBG�"1-֚XQPb��a�ė顜q
����ښ'�-gx{����`�SQ]�ι9��2�\�0
�]2O����#���$��E&��ȃ)��m��>Y(F�a�B��k�:�t��EԚ��F�	;k�a��ϲm�^��#jg;`��:A��J뺞����B#���
\}g�i�!�\s�M͝	�f�#����h��RI*B�����7+��#�	 g�Io�p�6~jdZi�D4�iJ�Wj�$�ք��\��F�*��x4�����#t�4��$���)4�5�@kc�{�V�ѣ���DwZEψ�2��	u�է�(q��S`�Vӿ9�|��s`�vD,���>��-���Y#���J%"ǌ�f������m�����p��F(��\��fn������ϳ�o�iK��;�6o�L��6�#ĩR��Q��Y�h\�]#�*B�V�/�?u�3�d��+&�]Ȥ�1���`�I�UH�&���2����.ɇڤ9��M C��I�f�i,���G|6�}���
f�/	�WP����B����W��~�G�D����VJ��ahL�k���)�:�d�EK0�4,���ڊӧ�r@��DV��fIZ�C��U�tGN�w�-iڝk�\X�[���F�iy����
$
{^>�p�
�m+�h¿|DHys!	�{��C��U"�Vܛ�S/����O�q�T�Zr���J�H/�(��e tV�\�}�@8�x��Y�D�{$��'�C
���+Վ.�xH�SަZ_�
��o��Ι�E��Lѐ\�1\�_yuT*�>�BY�����rմ�L1&z4Ro8�v1��+�"�L�~]��X������ \}���q����,
�N�+)�5Z@m�Z������ѻk�e\�r1��B4S��p���Y��O!�tx�z6�b��ٟm��GN�l��d��o�!T�� t�Sʁ޹��L�:x��7ble��>M&�k��z��}.�9�ؙ�$#���M�9_����BӪ�;D#ç����tz�b_Z��"��@�˛�����Є�y�H_V���#�%Y�-���TSuɎ��fY��`�b)�� ��aր�@�����gQ*
wWx�ĞrOH�v�=���ER3�t�ZX���r�����\��C������f=�����)<1�)��ep�;G;O� >��Z�+
=-�ycL0��p�)�$.x�z�/��x��߯�sY41�=���j	���9$<�N�"�N/�;Z�,�@;}�ycqT�3��+�M���	m�9_(Qp���#�J1#AL����G?j�nՏ���1�M�"�ħb�{Aޏ#u�V�j��2�Ջ@Z-�!W��λ֫�� �ZB'���Ky�8�@��Hx��cC@��zy�c���hMZ�m�P��f9��V�^B��Ҝ�'����X�u�~�⤧X��/��&?f�HP\�LU\gzgY��?�苙����S�7׍��SKB!�%�`�2��ba��W�zɅ=����g�É^��Crt�K(��\��`��>P�˂:,�1�¾-B?�Yv^}����=�b��>Q�������a�eR�FZ������B򤵕�^G�"١Q�*p���(P�Z�V1Z��+�eb���3�*s���z�k";�BM��͇f6�z�+i���ۋ�x�ӸuO >F<
�'������c]k����S*[y_:v����C�^�g(4��l_�B(j_�!6��(��;7������Ǝ	˿��m����ݫ%��($�^M�"�{��8���# (�2Y�@	o^/{;�(�H�f(�0 f�U��k���ߗH'��ޜ[���N��6�3)����U��������E��%�������t�e�=���C��D-�bq���Ĉ�'֬a�֪�����@�{ ��UK�=���\�Oj���D�P`3K~��UO:N��C����"8CK��3ȲG�	���w�,t�&�4��z��s�>��M�-��ގSy���S�������=��)P�Lp�1��m��3 �I7���F��"�4���fh�����o<1t�B�"����+)��~�����F
@����B�sUqvQ�k�����?.�i�{��[�Q-�ȭ�n�ӼO���!�|J������-���(�x��"�/p���8�C�C�e�vz'�2Όe���ŷ�<���2H�um��J"V�m3�!��Pg�DZ�ﭱո��E��s�3__�H�m#��p\�������t⽬�_c����j�x[�X�~���y�C���<�|N��Q�l
�8��--\�'�}�<;]E�:�H�Q�������tP.�} :�^f$�H7;�	'�֨�G+�c�UQ�D�÷��y�
�<�J�1e0E?�K�Z{�-�
(,�E�"i�jo�i�ą}�R��_ydq��W��a���:���|��B��ťEO}تն��R�¡�a��r���H/�v<_ȶ� -�!"�%�g�".w��'wϼߖ�F�|t/Ls�F���0���	㣨E�"�f�2	w==-V^��j�K�ep��E0ٌKYTք$�{���%�	/!
 1�����{��D��P����鞬��P�CQr�]UD���3P��U���tn_M�;��)��݂B��F��NMD�V�k\�i���;^��l�\���ݙ��2���~��}�&���O����-S��9liź�_n�K�Ġ�I�&�>���8��elC��Ң���;�Y����k\ץч��/��bG���ߍ�iT�҈�b��_j$}��i�[�6ڦ�)w��yA�hc�ZĀmm� ���_�س�72|��ut����o+3c�y_�	\�lߞ�ض6I{-A4ܳ���y�����+L?��oNt��`*��D�
黬�%��ŉ�=�?��
�_D�%U3I��A�E���7+���KB.X1��5��Dƍ����������@�N�L6Ph�Fl��h�^˓� �d�^4<�twL��ĉ������
�Ά�~��D�KVrr2��%��1��O}-�;��!��=S�2� �EK���c���#�܌_o\?)-�C�[+L�.�e�D��}�r�6�i��U���\���JM�,���)���Ke��L���@{\�If�H�ޫo�TP)�a�DG���+o�Qb����t�C��X��ڒ��˨�)�|0{�)�Ǵ�F��"�yzt^s>#Ĭ�B���O`�<�,S�* '[±oM�%���R�6�7���`�_�FB�~YK�̯,�	h���|�N&$ЫF�&n����;1z � SPr��/V5�nz���IaȌ��UH0ԃs�V2��_�����x�*#%��0�JnEۛ�=��F�yW럩��4hؿ; 0�ʐyr�/v��v]d��aM��擋�ML���u�<���ӥ�����<2~��1�V�D�`@���<6�3�m)s�iČk2�c��+�aA��E�,̉�&��k��򝬁R�қ`H�a`�|�zh���#v�'�o,��v�������@�����rM�PZ�3�
�riX]F��Z
���q1ɲ����B��sGt)��n<�����Ii����ɯu#��+�k]P� N�p�*�".�Q7��]�2�o@�vt)u��r��iʑ�1���/S�pLU�Ϧ��m����~�-j�3��$�ȑ���x-�@m�9`7��L)����ZЙ=�g�q�l�I�F���mx�Σ��� ׯ������%~����x��=�n�s��[3q2�a���̬���&���~kSkt���VQ��Z@�la.٥�l�;�͓������:��}>�e-��@#;�/��G�M=bR�Љ�t��"�k2
D^9-?��c�5r�ρe9j;,����?��"R����"2PJ|M��3}�h�K��/Q��FW�g�����.�1��5�y���c�P�L2,!�,J>�� \�_lp��,�O�6��K<������41�������-5Y�ÖK@/�y������-�L�nh�o���V�Bj�RqD����.���o�����a*k2�v6���˓���]��D��NyIL;Sݧ)��j���K�=A&�Ho� �Ew��f%e�L�SRt�'T�H���I��тY�ZW�S�����S�V^�$O��pZ�5���k!�Y!��Y%�Gll�	�(�[�@j��#*xݍ�٢J�dr	�"њ�%����i�y�_&��5K�֦�č��Ǣ5p�^vn\&p����_E����enI�t�[��v�x�O
&��Um�[-8}DR�b��1�;>O���҇��)'�LSnyK�-�@ߨo0jyX?π���P
�Ŏ۾:�<��t��/�}��U|�e���]�#Dץ�~>X��3�گ7�/eG�-�2b�ݷ���5Gh1�ڎ�#xj^��!ҷ,FR+��m����WyP*f��d=91�H�����;�>0��&g�؋ݦ����'����t�u��Y�࿢6���fS���T�?�	"F�����t�T�&�4u'�|��n�Τ�Oڞ�?��9_��|{���=�quh�`{�����D���ݝ~U�\�>�r�nIl+Q���+�[jC��5�������W�7E��>��m;&Q��4�J�t]��#K�$>4���2%eX8f��S��z@<�'���d3�P:c�����³�Q��Wn&��0.���f��B��P�**ò>��{c��4������,��|�P��J�]�2Wvi^}�o�vz�~�
{��$��t��T3 В�j���&iE���P�e����<O$Xn_,�=�y�s�ќ��)C@ޔ()T#s�@,b��K� l�B?+2��ჾ���+�Jċs���Cr=5 JsǦ�ݜ[���Gt8 x;@e�R�Hu��p@H� �&/��byi��w�si.kY�,��P*�Đ��_�/�pQPއ S�,���޲y�=�E��?(�["��D�2>�k�����~ԓ䄘���b�1/b�c.��s�E�2ˆK�8U���="��d=�p	�{���)	W�[7���9�Es�N���BCÄ
�}gR��pߐl:��0A���p1���Zl�?�A6�!�}�ײ\ے^���J���r���uŌz�/�����m�R��[��L+��H�nzOW8]b<RNƕ+|_h�g��� �|�'1� ?E\�:�*�ԫ�|V�[��5M��P��Ob4F��a۔]�ܤ�	�t~aq1�\g���n̈�d��ہ�P|�+� X�>�X�v���`��2����V�=�`A;iw���ü>k|U�$n��*�DC���V��plUc5. b\t�{"+�������J��'@�!��)f���[*#�����)>ɕ8`�[<ԅ��7�&x�ߌj�a���cj ���/��#�<j��,��G��~_c�^Ĭ���S���L;�$Z�>�q�a٦t�:%g�/��qL�q3��V�N��es-���6@�9�v�����8��k9�^������������{²l���W#�졓��dE�\+�����wH���x�^�&�Mxŕ��PFo;����EY�u�ɍ��֕���-8� �C8*.�Si����N�0M�|U���?��[��WGj�f����LH�^��\1�	C�r̄:��v��,O�Q�y9$��l�;e;��GU{H�!�,��ę=��������h��gҮP/}OȜ!�`h��aNb?@��i���i
�OZ�XU���g1Z�ZS���%�|���Ѻ��_
�D}�h��'V@��_�W�DhazD���&)��(��㊃̅��Ri��.ف��#�i�F�N�EE]��iw,��e
�i�hU���aM�9��
��w�M��q�*"�)��x��W(�����M�i˂�N�R20�L�'*x
H��&&Bg��)�>�9�"���	ϓ��	�ĝw��\�v`����Eb(�!��;hn��p{�a�l���WFi��P��#��u�r幖�[S�BT������a׶bb�\B��醴w�8m��5�����'Åz�-�3�&��.?£�xKd���0$FY�e��h��U)��-�Pi�(}x2��[��1K���mC˸�rpCw�ӣŐ�x����Z�n�Y��[��m� ޖ�!C]1U�G�L@Ct�y>ڜ.�y�j` �΢�LmØ���#	ߦ(�km�nƟ��**�<��Eu8��*ޟ���k�Z���NhVz 	�J��ge�q�[d��6�k�q�%8��[*���W��������f��rO�i�~�h����d����θ����A��uNS���:�O�?����ĸ��͆�߄�����`�=[���d�� IiAS�$��<Q���)Q�|�������=����p��5�Bh �.�/;b���DD�/����Y']��l,$��
;����&&��Jzjy'�ec�ж�t�T^�E�)�A)�v�H����s���q
�e]f�ɛ
1:dm/�|G�uOp�м�"vQ�A��\YTn�J����|(sub����#?���q��$f��'�,y?�K��7���Gs<Xs!6��r�֮p����H���������2��E�����MJV���T���	(�l�s�gƓKs���Y�Ao�>>��0ax�l��1.�.ǀ�m�'49x�ځ*x�Jt-��O�U��e����Gr��6*#ͱfB� l,#]�Ό��;��Ic6�O/��A}��*E�pI�=0��A����ycZW�2�I$�<��l��540�n�no�g���ŋ��uS���6<��y4QG�m�C\�d�R\
�haҽ��ԟu���7�e6���h%�����U�@O�-���5$O�
M>(.w֭jlO��Z&[�Ok�j�b�(j�tg��ybUgLD��ʺ��$��i0�n��X�Pjj�ǆ�EtI�?��R@��v��k/`�p��N6�z���j�.��b�oZcf|����\u@�x���b�	q.m˝�r�T<%x8�4�]�X��Lsd��h�a�xM�R��J����9���!]��P�CoD{��C-����g�a[���:Ecjp�=Q1-;tt���&J��T�F���<;��ג��7l߮�@R>;��3�j�-�A6�s���5����J�0�BU��?Z�F)|2-�oOs��������+U��U?|�H��%��bj<�j�f��z����1xLw����K`���1�{����ޅF�H������l���"�y��p�Ո�k�Q�����(�Υ�,+�mA�ٜ���RbJ�وxӕ��ׯS�y�7h?�Q�h�����I�0n����a��Tm�%%F�&�@������s��qW]&���o�clCn�}�%���~n�1VvL���k��tE�:�P���´j����?�����l�P�A����kk��*��ڄZ/ŭ�eL�f�)��͗rb��9")˿m�����w� ��b=%��X'���r{c����7�C[\NP%��zA.p�!}���啦���(=/F��C�&� �?�7�����tM���7�>�4�u�TJ�1�Q�(zN�R� �OJ�/C6�� Z݊���':N�Ew�����B��&>�O�V�}-+4�"�L�^݋X?�\=��ҧ�sw`�G�v��	�]N��uf� ���d� E�c^kɭ〢�*��C�wk�Gd�;�Q�V�5�~1E�"e���|�4�m�����ڣ��{�OzX֏N�Z�[��+o�u�<& ��u���sOQ���T>�X;{��Y�� ҇�{�ٴ�n�4��w�|�#�ϴe��Ox�:Y�YEP��ΠS�f�h[�����:Ͳ��t���:�{+��GSvKΐ�Y:�Oa�RMs��U鷣�> ]{��.�B�|���ƹ�9��߀,]I���Y�>�e�;K|#�!6_Ex�&Ug��x@1�i���27�Y�P�|k�5�%����(����K�Be�L��1e�X���j~���P����9��*<�+?4{���ZP�������&{6&�N&�Z�)L������T�$�FY�0�6
�����_f����a�q��0Q�k���z����|�8a^�aB]�X��j <�>5')*uA1�_�[k����ԙ�\�I��'6;��3~z��(�>�*�qw�{D��{�~m�NN!��,�]rP�،i>���g�o��ίK�^�JD�)�A��a�,n����0Ib��MX������:�J�hR��ؐ�=�� �$dK��i9s?6��}��]?M#E����k	�������?[K��dR�c���eW���\7����x�^h�O�ÌT���C\+��\�~8�c2�hx$�/hħ�r0�t��`F�d�8�۱e`����+,���j�6�M�w��s�ozJ�vksz,�}���	�2��X�!���5����0s�}�R����G���,hvMM����_وg��S�o�!��M
[�f
���OJIeg�TR6u�+�sA��-<%���M��?ǫ�e�<v�~E`w<3G'��'D0<��V~�c�7�Ю���pIM�l�m�p9��Q�/\�JT����9�洧�*��m���͉�w�pJі&ժ��U��J�p�ȁs���z=�x�=��T���Q����=z[!�l�:Z���d�8]a]SoN� �(Q�X*��J��	���zq�x{M֯�t`��(���	��yCn�$R�a��#�SR�(%���K��ڠ[���+��1!�Bf�?�b����p��!���o�W���S���7Yv����0?<�]��n2g}��4�	�X��1�J}������KY�$�m+��5JR9ܿfS>�N*Dӎ¿��r��%���ߜxK�Xy��!����e�g��BM���DU<�4�b��� F��u���d�{v��l����i��D�Z�W]MrXc�wb�=v�A��g����A��]���V����D�M�i�Y�H��Zv���+Y�K:��P��AZ�.������� ��Z����!����`��ɑ�!S�B���w̢5�\�^Z��d�ZwE1��y>ZTl,*l��=z�߇�'�R�@�l��DE���[���B¿������/�=}�/.uE�CG�&'������8N���,�������9�>z��8I���T|��IJ=@1̜���߾vr��|��`��T���?"�VY� K+���h����f�SD�v��siĆn��+ e��+}�m^"V-z&m�t�.��@��v�詭"���z�'���M�	6Sm`C-����}���A�~O����+�a�n��T��>c��-��\-�Z͉6��S��1��;4��﨑���l<hqsڮr�V"G��n�M�q�<D|l���Li�Y��O]B1��K��hR�	0��H�W�N)G� &��c�[�4�Y<#h�o��k��ds����3Ic�?��g3�}��C��4�5%+�|���8@�i�}0Ӎ�#>���4)�P�����!ہ�sn��������51�*�Ƕr�Ɖ"�9�E\�]�M@	>G�%v�~6�;�{�����BMmЪdZ�g��ӷ�]w��+�?$� �A6�JxC���f��{l��xr�V	$g�WU�XRQB쪮��\�0ڊ������;Rk�4�f�����x��|������D�РIӑ#������5jD�Yqn�P٨�c��Z�#q�.J�x��(���^j'Ю��09���s���K§���b^	R���-��-�%	�%�J��7��Q}Z\E��/��:��Π���J]6�oy�9���o`�H¾ ��)�빡m�/�߹3T�>@y�Q�1�����Bc2_��e��/�z�����e:g�����xI�ȹ��$�Pj�e�X�i�{� ���6�TL0�%�:Y��U���s���oI�N���,H&F��/ �ht�?��k
��%+=Pt����rcv푋ͼ�Q4ɤv��P��S(ll�k�I�/#������|N����x�h�9V�>�b��c�S&]~�GR$���eH���8j�?�\#�i�gnZ,����]��6�N��/`�p63EH���$[��.�����M�.��n(_+`E��x�8>��Ub"�@��ZS�+ז�4i-��HX��B�!�AG�� l��
]�	O�Ȭ15�v�g=�E)����'5:ء���K4���/��r�7N`QCH�"K#LVaRFa�W���邺p�� �T<ڪ��ل�~%�Ds�c]�JӊQ��*%5�
�Y0[�s�Tc�ȃ��)h4 v�ǚ��hI��1��}�ht1�
pa*8N�|ɀ;��c28(�}`��^C��ɠ��/I�G�@]:	'zN����/+��M���ft҈x⦹Q{n��W�7���"�iW��U��/�c�!�$��i_숁�h5l��m���ys�V���JkFd����[�[O�$�'/D 
�g�:!sT��eӖ.��_��o�D>f��t��d��[1���٣�l4����v+�`���d�*����a["t_��[�р5:��.��;��p�^����ߊ�����ݙ��ė��WS���c�s�o��:��m+�W|��!D�Ų�2�O��E��?"9�� �?s]�8LLZ�t�?�{�#�>�C�`+���7r�j���%�[8x��x^���$Ę�'��9ќxG3���s���sD�{�w�nV:FQ:�i�(�:�Eqd��~/�/$N��K;ӻ��;" ��e��z�^�~XF6�7K	��9�>f4F���u�qD��,h���Փ��x���z��4�n��f��}ظ�C�XsU􄹊o�}�I�@�i@i�o�k#`�t���Մ�cJ����58�08#/,mto7�`��Ҽ�V�-	��ߢ��1| ��ĆL�a����,+�h.V�H����\���%��� �b���uG�����
[�o�qt$����e=��UC�Ǔ�*g����U����>#Y%��?���4������Km�w�M�X��u�.��Q>V�*]%��d����KzR7Uޤ�?1=n��?֐���r��Voh��+����#.T�e�V���W��.�CU��[�(�3[��V��S�OD��NO�'�'�]h�:[�V�/f2�L����i��IA����
1y��f,[� 5�_�8������5�f��X�"SF�!m�9:0��n��ɉ�tz�̮J��o>�~X��c�)̚�0(r��1�bݢD�Wp�%��E�:�m����j�O���	�M��W�8%ud5
#<I]���[d�&�ƶq]%�6,�긌2�DEQ,��m:���D��TK��G�\�f�ʗ��D�Ct�U���q������#@�_�V d�yxg��X:5����'1��;�ҵ�.�w� �š7�0E'l&�o���'e
�+f��c6�썁o�j�gJ{DB��,�'X��n��"��Ʈ���`pO�T���������ˢ��4�;��7yRL�ޜ�,�[�y.:@r@��_qa��A66�`�~<=��l>�ֳ�A�t�֒�6?����{�m`3uz^J�:���Ɂ8e6U�x^w,���F�f�QXe�L�|vH�#b��r�C;�&����D��T�=Λg��� ���@�ߒ��3X>�R�K*���*��w�g�C ����2f:��,?d��͓���f٠��P~n���V��սs�V�|~l/�����G�v
.�y��Z6+tl�b7ⓤ?�0��>T�@���o�O;&�zkK6]������-8���ye��97�	�1{!h��:\�#M��������hh@tM�yB�&�	��3�I�cx����� �id["���ܲ5V*-wp67��n`��a�A^1I	M���9@�t�+���\������G��*h���%F�&E)����5]^��I:�v��X�.$��a�"ğ����f�a�c��*�^W}O���<z��겁�����*v7��%@��8����Sņj�
z����_��JFQ��ݔ�-e�Db�a�߿e���Uu5�0���㇕��$w6�NNmag�F��@8
��6��(>��2��qlc;���$T[��O�\�6->@9���Gt�u���A�'Q`��"J����J�����N�'��o3
�<>�����i�+�h��Ps@�m��r+�[鐡nѧR��������^$8~ȝ�F��s��[�tࠍm�?>��z��xUPS�Y�9	j�Sai�@��d�&d��mc^]��.�!��l�);���?����dBݽ�~��~��qEi�;�{Ȉ.�(��g1)���h����T����<�-�Sm�k~~�aG�\ķ7/�U����A*��|����������H>�+��򉄿s��i���ПϨ���pl�y����>3�N!�hX����o]��7�hA�-��7ߦ�Ux-����sF�N����峲ﰛ��`��[UIY�t΍L`�	�N�"*M*��f�h���g�^����Pt��������W�M��y�]AwW{PoN��9�TΎ�Jֲ�����Yt��*2�ꌈFV�B�����(���QM�@�C�k�ea�}`�,�3��/��r�����\�;���kZ�:�������uHb� &��|Idp�s�H��(7�1]x��bd�H[�����",?n0�}5;��D��Cޏy���pm�Ƿ�N�L�;�c?=|�J�?�?��y�K���b�IO �hh���2ӌ!lۣ@��ɲ����M�j��qM����sn��i����z�S�Fg)�GI�B:F���z�:٬��M�U7g�IS��
57��OцnK��n�Bא�&-�KLf&���a8Xa��*��⋽ ������u������� bl��[�#�Nl_��#�����9@��l���)�w�㢉��U�=����ҡn��_:�t[ي;�j�z�V-�PY����M璶�����q���f�z�.�6I%����i�j>�p����\�ZsM�λ� ��f>+�h��K�1'�ڧ)\�)Όk�9�m�~&��=T�&�P@�1�Io��A]���4��sh'����Cz<�CkcI���B�Pq����Q��������T��쪮���tV��;��({ܪ��7���S�����w���g�?�K�E�&J$�!�������+��563/���nao+(�����T(�#�*�����?tߑ�U���A9�D\���4�n���[����m�����:AE�H��O݂���P`t1w�r���P�>�RJ�̑T���T�:�}��Asm���Q׵��/R�Ӝ��*��d�+�ۋ���|T
���B���I�n���2�uX���v	�5���v�=�u�&�r0y;�Wv�����,:۶ژ�� ������C�u���zX�O�Ҹ@�`��d	:sU���F[���S1��"�2���n��u3�`�Y�6����3�aG�����(��*�X���jw�t'vB���-ls��5,c�;:ط��L3���X���wazc��� ?�R�n�ʷ��)^�!��������亻
�U���Wp
�=f=[E:l����!��5�_��1#?�v�&T�ۗG�Lk�z�_ܞ?���viB�w<L�S�4ޛ����,62�v<D��j��D[fIX��d��Iy�-p�O�4^ôjB< �-���>��S7��O�69�?`��X�ږ����/���J��vk��T�B�1��o7���T::!�-�B��b	,@6ײye����P��3�ntnz�<�{р]Z����]P	��!=U�	kQ���ط4���R���A��
����4T~�M�l1V�*b5� ���wP�B"���ϙ6B�e�%!������fW�h�U�߽�k��ȫ��I�u����i��c�M�������&��?}�����ŕ���7��[b#�Ͼ}n��Ԙ�-�L���,D=X]�$*�i4L�L5np��'t�ՙ�y
��H��r�ڳ ���K�B3��٥���Ł�V̔�c�8��kAU6- ��_�FA�oK�]����Csr�3�)m�p_��D[�� V/�'Ԡ�Wx'�nP:ߠ��G���.��3�w;������[j#Ν�%D���>��h�&/�v��CMx��?��'Tͨ��A|�%\�(~T�^6�zD�L��e�i�b��4F~�=f���jGZ4�g�]��F�ʹL������K�>m�/�V�`���-}e�s҇���rsw�P�*��䈋�Ļ��A�P|�z亹�7�U"��A��8;h�m���a��ƴ#P_���v�?Mt��x~�QsQ�����Ik��5{�=UZ7��o;�n�-�ph���pB���w�0���lm|�5Y�������Z?��|w�Ʊ��n���:z����g(���u� �}��xG�(��C���n����bz&�1Y~����^�����$���w4n�e<͉�;Ӓم���t+%~��g�����X%H��"aA4��A3
������]%��
pT�-nq��j��ܼ��%o�"c�	�![������;���>�y��WY$L�_0��bWr�L0�� ie��^߮wf�����ㅵD)��XZ	���^�3�Q�+VK���/�5%�@e ��+>Of>���m���M����$��2�x����2��>lu(�.�{� �5�������y��/�.�z�eR���"����oY����$�]�P7~�A����]�.m��ڬ]
�y�qC��.��䈱�_�]���2�Q3r0�_blEn�w���2��^љ��S����	�M,Y*4P��%a�9W������t��п8�8Z�K��Y{ΪAz�m|�ajIszu�z����-��1�Ŕv��y��d�ƴAY"����ۥ��nWڐ�DY>N��I������5jf#Yg���g���^It�	�ۆ�@�9�%)J��P�F��*��9���f��o�vj��(^R�~�. %��AZ���o�.�Ah2�Ns�/21�>a���E�V����=�G�Y��'�^�?�Z|�� �3���(,�V^��j԰��;'�1�MqN @ؚ��6{�?�>x�_:�٪Q
c�c��3��� �.�N�GM6��L֤�AVݵ��"������0�`�Z����h>�TI��6�ޒ��_��:�k��׈5?���q����ud�+.^�J��o�:�ӵ'������UT�5G��f`ׁ��r�/���O��&�N��
ږ�4�c-� �U��_�±[�(�O	Dߤ�����i�U[�
o�uh���!�F8 =C�|0/D�;	yb��ɇ�23�����1W�K��W` -L�U�Ix��C#����ta���>T�c�� ���w�;�UtJ�,j��v1�Kq�.`#;�E�uԿz���sp�
/0��w�� ����ŝ)*��
tk)[����'�7�wgZ+Nd���k �@�t�Հ\�S�b@��#���	B�ķ���`� wVG�˖km�T�b�6�����$N�\|D0-�x�oD����0�y6u�)��m����l���cl�FQL����V;��w��a���T	l��_��H��8�����+?J�PCK�$��?��$�s�]]�G>W�l�NS\pr,:,kk~�#�Y�Ԝ��1�u�@RLT���k�c��Y����5������u]wxoF��o��C�2��8hX�K�PV#~ʊǐ��6��Tx�pX#�D�>��fUHS�ۿe ��0*�0��^�`���j.v��]D|��L�@�ݏ�Bʤ����Ѱ�b9"S������p��Y���uӽ�D��FQ���H�JBw���"0��ӰEȣ�Z�ӗȫ��N���,��B�ο��c1곚��g�*m�����ӗ��M� ��R�b]%��Y��E���~D�^�yP��%������&t[fD'>/���o��͂��!&�m�t��:r%V	��U�V�w8/{S����ߑ�,�lc�y����e����ica��aC��j��+ь���4��׀GC��K(ޫb<��7='4��1f���;�;t��e��;D�8��5өo5�X�,�G��Y�a5��%a.���{!�2�MǋM_�1������>Q�L:c���]H�����LD��;���}��'����	����k�Pp���|d����qۈ7��HwYia_�s������ ����8���P��2!џ>���'#����])n\
��G����7�W��9�c��H������/9���Jm�՝;Q0{������s���ev-m�O>T
տ�0^ivڹΧe�W8����%�ބ��w!+)�e�3V<�v���������p6A�=��c��|���ȳ�����h��&��+����@H���Z.n�k������٠�r0���}��r���ϝ��s���ҿK�z0d�R���~d�twc�ňx8,�E�n4�rp�j�u[�Q�t���4Ҝ��r�|VCQ���Z�ҋa���O��5�i; ��0�uu͉�V�l�yۥZ�`t[F�~*]k%7�0��r!W�gUcb��1*:R�9�yռA�Y���R�+St�ô��=F�K��+^���X�Ʌc�9!X�C�b�{�YZ_Ю�n�u��Q���u�5����;E3<����$�>_Tџ�{�3��=D��x����z�<sI󕏠��y����$�qg��Y���K0���r��:1��SK������{�waP�R0�)�<S�P�t��M@�8�c�w�i�*�� �t��ї ���Sl�- �Y���Lxϧ8�
Q�pj r�j�im��6�,��<4����D��C��T��$8m҂>)�D;�身d����xk.e���A�Ua6�i���3���H����8�Y���{щ�Շ�|�Thܔ�ʑ��@��u�Ƃ����>���SYb�n7��T�$Ϙ��`�@�M�R*φ\<�ޤ�_3T���l���/��$��i�6|H,;��T��@���e�l�����Ƿ��F��@�$����*8�fnN��8�dpb%TjjT��f�+\���/W�<���f�|Z�1^9#������������{�qD�G�n��[ng�"d%4���/twUW ʸ���!1����� h8�6B�ě{�F�����^;��{6�ɜ)�x��6��03�ӈ��"D�x�d8��G�72I9u��>��l]��}(�P������Kܕ�DP+j�ݑS��1�ח4w��UAv_3?"��6q"�$��d?��y��͇��lX�|9G(�Y/�$����1륃u`�Y�n��!�)\T�Ve�Q}<%ſ2�/���#Y8z!D%��L6s���D���P�8q�k��K��W �����s����wV�d�_j�y��"��;=���}�(W9�f}�(^�����m�gn�s��AOf�Թ�խ\=
-�P��<��4,�VP�O��r\�K�j�_I��K
ow*�a/8Gi�B��C���nY�U��K�;E����l����oSk�
qs�±�"�؁��H]���Ec_�*K��ZE"`�:r�j�&�|��Y\c���s�cZ�=�̰�򸷽��F|�:�;_�?ʯ�#$�5iekI�'�D���Xk�s:k]�+a0U}ΐ/}�YϤ���􀇺~ӝ~I`n�2L�ž�����������l��I�uf�zQ���&���2v���;�.�e3i_]5Tw�H�r���$�R\�Z�R�����&��!�.�H6 �iAs��u�#QJ�����4�É^w*R�*�E�V�yY��H��-��u\�rN�'h��L�(ʥ�n�AUZ/
��	�y��(W���	<����.��)�)�fT�|�l�+դ�!X�U�9}����d��j�2�� k��D��b8*�W>*pU��7��Z�Z{����|YD��k=Cl{RL��c��-�y��9F�h��w�\��~�#�{;}�{�|��ū�f��v٢��z��IC�VJ���J}h����g�E�B>��7O��F�e��!��~�?�:�bR��R�>h+�vuʹ5F��1��hxCH�:��������H���_Ik����'�r��������'Ԕ/ZDL��w�6�#Ö�R;ɡ3<��4	�Ut�~?�?�>6b���x�)� x�
��SY�/��w(��}
�]6dz朤̜����ǧ���!rr��,��Љ�6X��L�VW��Ne8w!"�?jye!� �J}�Q�u�ƶ�V&Ƙg�ٝ�k0Amg���o�i2�w@Zv��GSrA�]�ۢ�y}PZ�J��%�}<kl*�6�GES�}��g�L��?Y�/�&*(��H/qs���dJd�q�13͇H���6��w,����L{�p^bm�-d��d�W�7I����ܯ��m(��E���{}����6����鉄�]�k^\�Vy���M�!M]�Z��/�>R�A��-�\9��[&_->6 *S�����㔣	8!�Ć���'�'A,*ӝ_�{����%*l��!���s�Gun"gR��S1�43|Ӛ�`K�>|�t���Wc����wM���9���|�Jp�oܗ
K�<�k��3b��V�w2�©� ���v6�^�z��k��;���!�]� Ų7�4�i��_H}Eg�\�#<�V��z����/4��M��F���dm�pҬ�=ȶ���Żͯ��ő�$T�+�7;�
�V��&����3���)t��v�у"J�t�j��cGߛN;]H��1 ��0ra�����]�$>�4�.��ͷ��t)����������o������ʯd#��!|��yc؄D��M���=Vݼ�����`1e�Kp�E�o����7_�pEiR�;�%�Ŝ��/rW��)p��'+�HG�K�����>z�g����m��)�x`g����.Y˽��c�܄�:.3Ð@�IGu�Bi�3a�!�bPѻ3�@�9.��+!�`	;u��$��ya�q7�*U{��^j.��?.����`�����^:�k]�j��3%�m�����h:�zO�&z��ȥ�6E�:�I�f�rt��cG�7[�s�}o��� F���We������a���,:Ԩ	t5���/8!�
#��W��W<��T��5АE��$�	��:*x�b�D\ψ6��%G���z��b�;_B�7�s~Ÿ�?C���Ыx-V�O��V�Nh��h퀑��]#����3(X��2l^�Ԛ����"���t-~ �zi2w��"aq�H�Sa���\qnmV�o���(�[�����&e��Tf� %��UM�?U=Tlr�a=G��^���k��I�vģL����z��ձ�['h��9R&'����#;�@{��0�B+�}`��������M���<��'�m���Pڎ�T7��;�����EP� (�w�������fYn�V����Y��0�����y�!��JYg�U��
���ϻo���~ˆ͠�S6�Y�^x�ׂ �p�Y=���hc�WrL����w��H[�n*��_����qXھt�2v���[�mT�P�K_?Ʊ_�֋5�o��d��I�\�u���R94�$uTN=	���m�A�-��42u�þ2�������&ݭ�l�qBD��x�[f7��^���GN�t�#�ғ��s&|,�O�7��0LG'�W�-T�^�BV�Ӥ�ī���8��`|���`��~L��0��D�Ng߆��b����]�p07U��Hv�Gi�8-�hU��8��>YU7�	�^��	�A©V�����ȅT���h}z�˫g�՛��.���f�r�Lۛ�ɲ��4�"�2d�s�K�Ē���ʏ�-�1��<���p�r���t\��������NZ��p}��j������8ȟ�+��x $ܤ�"T��q�ފ�`F-C�	�s����3}5\Y�����9s�r���ޔ��ui~��3�t%1-B�UD��:n�}N��C����SY�
gϋ��Re�*tq1b��H�*�vu���������֊�N��g�N�};�lNc�4��>ޤ��,�1��b兦�BM��U����-���E��$�9q�@�D�'�$L3l-�x��!�c�ۃ�<�����P�a�|` �#�,<�VKh4�(Ȑ�@�g�d'�:,Z��]r�ܹr!圯%�&<�e,P=��v6L��?�����9$���7��'\���ڡ3��X&sV��j��P�Aj�d%nUur:Q�Ƭ��~�[EFq���QL�8)r?=������ݭ��y���\������%H^-�>�͇F1/�Sx��Q��Tn'���ù�*�;B��ϣ��dE9����`����`K��1|�t�/��c�8�Lm��Jm@^7��A��;4���/1!���b�ځ:�T�{cͧX1=J�i �Uָ|{��/Ed���o�gj-�z���]/�_��s��Nd���
��Lv>��Ƴ�"��Z��E��?�XH�3P	蜽˃���w��	�q�T���
�6B�����.�����=KPK�3nL�`�>�K�j-!52�+zY���s�]�tR$��H�C�~�M�o⦡��	�ݱj߸ϓB
ʑ����x�Œ����D�A`C�vsp5~��`�]YC��L��V\��q�.��)�^`���)��LD���1l�E� �j�t��U�U�D�k��\�7T�1�� '�����o�b�A�Rէ�0'!�G�i	�fz�X�g���s�q$?�M���"ꝩGU�&����X�>�rsj���G*�%v��r��" _���\�u[>�T�Z����`�0�?J�t�C����)�g��6�@Xe��N��)e���{�J�GE�j1"�����h��a������G	�l�	x�pE��P���qֽJ�w�dY��ap�)�R��l�&��ren�o.Zm7��oа�$_���v����Z�jpq�\ʝ���+j�é�u�����w���>�*A׶+��6&,��� ��j�7+�.��@��g��TǢ��-��a+��#/m�LnEZ��&Y��Z?�]�p���
���7��6���^c�P�D�TOlT��9�E�:]�
D�k$�{��w�;>����NWGX�~ua�w��3���O5מ�^�RhE}�S?T��#pd$XE�!E�� ű���u�Α�8��K	M#Q�jzQk�����zs��8���������v���L���s�$$r��|x�q��&�cyZ�MgT(��t@����"3�>���Y���*���&��+�����#8Ț���\�G�=�k�7˚|8�Ÿ�.���V�Qz��rK�U�|��������C��;`�݅��}�mKd�[a��#��2�6%@
1��U�g����ֱˁl�%�g�>|aH�FaY��WSk������r���v�W�#�ہ��*t�g��k�+{2�!Sl�ĚvmO2!7��� 3���ȏ�hzQR�,��r}��g]��m��b/�a���@|=۠��0[^�brJ�,Y�u4*�-�a �G]��6�M�0�"]LӞ����e����������,���Ņ+��X�}|"��f�l�P.�()S�[ٕ!��|��k qj�45�?"�ܷ��hV65�F����Zd�Y8=<t�b�	
[2�0��u��L��Z��[Za��``��i}��U.tf�9�4�<�1��O�0v�c��a�m;��b�mx��������d���  ��q'Ĵ��&H�ōE+gTչ�%���\��ΡM7$��.D��gF.��� �i����[N���t�H�'Fm�Ԯ̱�,c�Yv��d�W�-r�B�y�����B�$<�\�5��r�Ռ�i�QG5���@��pC����l�_����M�7ۙ�t)�q�^Aۊ��i����aJ����W�"��B���Y�5>L�p`d����qB9A\��*u�>J(�F�ihl��P+f���ڈ�H\�~=��A��zcf6��^.����C��ʓ!�>l�łut���Y���E�R�����j1�d=�$ɡV����9@\��R��e.}}����lϓ���S���]BYc�(�h� ��`��'��z�rhM�Ԫ��x��`�X£@�����D�)�ߓ�p��4Q>�䣩0�̚�=H�sWC>M���c�}i^�P��4=mkSG�p�R�� Z񫟦�`z�L�<��{�߃,w[�:ܺ��{]dSP85C~f^��[�^��O;��
p
7����@���(3l7l��������$-�C�MW=�I��iiǘ��F�o� \7�M���TQh*(�<�
��� ��:� ��}���]�5x[w���㞞9yu��{���V.郪��:�Ț=�L�@�`&]����Č+=6���k�w�?���l� ��)�7�RW~^�_�g��n�D%6�ζ�t8@��m����o��>��pXP�v��{%�|9)d���9=uQk��z�`4�
v�-��i�,9%��'�*	�X\���=+����$�yZf��t�C��������%�ˀ��ꞅ��xg�g}xȶ3ۿ�a���;Mߝ���%��_��)�9ۧ�?�T}T��al�җ�l@��f�䁿�%��8J��N�z�h�l���w�	�	R{	;�V�H@:A��(�j�P�7������
��w�Ut�b~�QgHdq�>y��)R�*���nʍ�-n�VQ��e�u��viy���Ó�{���aV����h��kB��y3w�@�
<���-)��&a��fua�u���bE�rK�-�4<��*Y�����_�[�h�������
������V���?�R�]ڷ�-��b��+ ��aBow��=e<1|�u!g5%��Htm<�������j������o�e&�;$șh@ �P�Cw2�<�`��9�Z�n�w5`����=�0�n�Z�3RZ������r�~BŊ-e�е)#�q��#\X��.��}��&9�G�E����׎g�A�3���H�l�r: i0S28�����7mz>����b�Cof�U#�0`��?J@� �8�����	�Ⱦ�B�
�b�u~ >,o��	u\���*v�9�nPm9<���e���H�x�$v�;�]����[�M��k� �jk����|� h���P�8���KA�,��D�,_���b��2���@q���̶{�o��DG�����������[���F#8�э.)p�}oW��ᙾ��CR��
���qż������M��x����spY0ŷ.@�P=Ȍ|�b(8�cK�$�cgμ�Dh��)ԗ���%&;�6�d���>��|E��bO�">@N�\ZA����G<e���h�F��(n�ZU؋}x�'��P��ʟFvj�^喚a��˓8������9�&�i�_���j��7�8�O$�	�T �$����]#�~B	���mz�vw5�VbꚄr�4½u�Q�mFk���{��x���[~bUh"�Gb`��@�	{|2��3?V�Z�u�D�Ц�m���}��öu��.
99f��ʼh�e�짍b�A�iIX�8i4>"���x����U�����W�xw=�m���kw�m�B���1<�+�_���S��h*�c��Ikȵ�'Q�&f��<2���cT�+�}�k�*�d�
�:�nPCsN��(G_N��,�[(��kc��7EY�́�}�Tәww��ZG���}b���eG�\),'<��"L�D,C�X���cXf��'����c���ޒ��5s���S`d�G6���}s�a�Q+����	9$K/vIo�z߭穁O#��y��)���/���*S{��o�" -��	��so��U�����l��1e�&�1��&��$b�9|�IB[8�7�`�A5�J���C�I�P���ڵ	�E�NeΆf�+$�o���i3��"��6pSj���$�%�X�Y�T��zk>V��f*�C���)����u�7Ji� ����f�t$t-�K���~���,#%MJa�?�,1l���l�3q�j:�i��!v�-�_:�у��+L�dzy�X�h]��S5�ذ����"�`���W�E6*��!ϳT�᫙��yi���Bԓ�A �%Gt��cO:����//U�g�$+z����e���r�i1l�I � )4�&:��=�8Hd2r�Qj�D��pm��LID�$#���.�5���),�Z��o*?�Kk�$���h���;����oDd�w��gM��7T�'+;W���懥��0o_�fř��x���ܤJ���D���tҕ���a�E�_�e����,�%"	6F�VhO$��)qa
�q�ʓi�X]���� V��O�[t�9i9.��aD���,�7E�0MF�}���xƗ�m��U"5�a�Dw!�'��yZ��q�:��
�%ې�	Ry�����*��qǶ����>� c�/��0-�N�A׎�	i��ؤa�B]�H��	��awůa�cE���F�U�\'Hh��h����]�
�2z,8#���)F���y��q$�����o�j�{N�UVǗL͏I�Y;�����sށ�/V��i��JeF��]B\���Lv���B������^Bd��$���J�L�s�D�����Ч+��Lv�箩C� C *�U�'�[��+�rsװ?����x�����Pϛ��ﾴdB6H�/����J�*��(Ʋ�I�K���g}�b"wh�P���� V�<D]�Ή��]E�Κ�����+-���y�'�BS���� M�����o3���9���1��<�2I�#�R��O��Z��s"�e�g���U<�}?���h0o�{��mSj#t~�l����Q�����ѿ��h�v�=���qq�������u�j�m�����!���6��
;\�)�8'â���w���Ü�E!���J����$
����:��Ż���G �-��`���$�5=�A�tp�,z-���mc��#��-��
���㬋��'�Ǡ�֭�F�K݃�T�{i��0E���|%aW!bKބ2h��?0L�aC�����JC�u5�z�+�(���� x���M$u��PO"�<2?:d7D�ؒ!��/����6�b̙I�d��]�,Y|��I��|����I�{\�7'/GZo���w���RM(3���qKŤo8/쌜�+��oz|cҚ��:y}���4ET/zQ@��?���S�$���������J�h+��.5r����z:�P"�Q��V�U/Jd�c��j�J�CLVQZ!KP�F���W�iS�p2����CE,���Z�<j�oB t%<�&R���*����~��х�(�ن�����{�����������y�;2��f��?���}so��Ҡu���#��n��{:�*�f�[��Z� q����y��*Ifm��/�.N>g��=���"	c�k/f/5��R�N��f�>oۖHH��
���r9�g��w�����=��o8��@cCcM,/6M��������-�
���DH���"{��B���7�cO�l�m	P�n�1\KT�4��e���3Ĳg�\"���
�c�O�8cJt�q$�1��h�7)(q�۽�7;B�?}��<x�����Qs�����G>v_���ƒ�g��}W�l�;��I��~����뚔�^|m���[�Ϫ ͭ &�P�R����'�H��9�f����$�F�<:�,��d��^&0�cqg���V���� I;��-�}�&MJ7���NH]P n��o�A��w䠲��.{��Q(.�T%���&I}/�x1wU���]�e��l�r#�st�HMSi�5J�݂��!\U�A��ن�䴛�W�7�_)��3W��1��w����z��7ԠsŻ���2nN�9n4�ST��3�HFM�qKP�2+p��ZG�T��n�k`7;~kнJ��h��(f�uTU��?)�^]M(g�%�=C;>B-����u���6/�uQ���~q�}���>��	�R�O�8*@�>�E?����jc�Z��%�AV�=Я��5�إ����tl(-���8�+�ĎRm�O�>I�U�� `�<(�����-z�f�}-8�%�S#L{O������Tr��3H��t�3c����D�7!��p�`*�h����ن_�b�g�w�q�����*0օ�=����+7�L\@��2	���'�1��͡�"՞3��p�����]%$��-u���mw4�K��YhP���=����.� ��Ձ�R��Xb�TC����&Hݴ��Y�_2X[��y����<�;N8�|PJ���TM�&0,\���}��)dΚ����(�a����>%��yܛ��TU���n�,J���}��_����N�����!�W@�|�	�N��.�#���g��ǝph]�Uj��FC/����׋!ϱ����\�'�E���
w�A�chC�vJ"��Ֆ2K��=��x�BEYvH�)g	_D�Y_�C^�х}�}K���tt<J�6��2��Wt%|XW�J�7��Wʴ�n���}�XD�
�~$�v�3kS���q�a�����_>��wY��+�������˰P�8�9�"V�[���ι��|�A+���	�av��M	d}Ź�T��C_���Vq�:�M�I��-?��w��!���34o3�*|�iS����:G&�#(��Tzg.%?a�tJ}�����\�}�Pp���9�
t�-&�����|躻�8Sd���A�`�n�����J��J�$��x��z���Ix�)��3�5ߎ����O�̴Vr k&�G,S�)C�f?Gv��v�@�d�Yꢩ9t��Fǩc,�%�1�I/S%wV�0I�MH�]�k㉔B(��Q��iY�q8�e��0�;�T���^֛�$�c���$�W���߃�q0�k�g��g  G?�r&�gdUe��m��T��Y����'�9h8�*1�/�����_V#�kJ�2�����b�����@�PJ�y��P|��V�rJ�X�H4��hT�e��?�����1�v~a�8�`�>3� 4����D��ֵNI�
�%@t1J�Y�fQj�a�_sdk��J�z�O�#Qj@C�d�b�m�/5�N
��
+V��8�A��$����ctb�����]��3|8Qp���i� 4�nG2O� ��,ʭJ��n}3 �)���'�1E�$�퀈6��J��O���M���%���=D#|be���-����4-kH�~hZ<�.�k����d�R�6���f�LE O�z4��>�'���n�U�`�bG�SJ�n��6�}/���qҚ/��1�I.{]	hc�o��t-ٍYH2T8����frCR�� ���8�SW��.03p}']�M��˸v`4!�j��F;�V��_���ă��4��a��1���Xi	����T��Ju�wbU�,lƋ�z��a$�+N��z��� �`�$������~��'��,VjZMJdͻ���� 2��'�~���ͪ��p�����8����)Gp.PI�k�,�~�
����������Y3���
���N�Z�@��]S'\�`˸����*�קL}~��i���y��"�=Y�jY����8YL(��y�ih��%����22��N�_샧��ԁT���F��""w�b���+1�^���L^ǻE��4f�dsZ�Ƣ�!����oDK�-gRm�/�t���{���PvLj�;;�I��*ۅ��R{�,7c<ή�{�Ρ�\WY��폤ˬ}>I���:��2$��g3�c��j��u\��x�����E�ۯ�{��+ز���]��`G����"�N�������������K�]P8�q6��F�蜋>n�� /`q��4K�"(�Ns� >��F�cQ�k�9.V�b$��E�B곺�%�����005^H=Ť��ˤ;��Q'��a��}>�[��mF������M�`��Վރ����XRj�=S%)w!��=�5�׿Ԗ]�)��m��C��Ơ>���:�/�1�7G��V	��7[*7q��F ��P\�m��3u�/��X�/�ֽE�'�`���_$��߿ C�~�A?�$c���5�wG�W>�V:�?b���UE8�KR�q�HebV��1���f��b,7�
�4l����yVS� �
��v��-G��&�0(NQ1�J�'�D���[���E}���j�&Cv&��ɰ���]z�v��*|��4��Es6�P��BKg��]g��n�r�ô8?mN�$�� ���1s�GЊ�l�����p���c���y��%]懺w�%p|��d�_���x��t<��:���ٟIYv�ed7�4��p�e�2x}������Ke��0Q9�4�����l��:#�u�E�Y=��(I��"{�fE��V�^N��GN�x�/n��ّ�@�����RL���h.�����V諓�J#T/8�Foݪ��2hܮ�	Y�J½�70x�ثPZ��k�R���L��l	+]�����.Q��Z�-%�5�%��Z���4�����O=����BR�"!A�\��G��4�K��b]�%�ů���sK� �v�d̠�~��z�<Fr/�����6X�-ٍ��x���<��U�`&\,Ɔ�j>��ݦv`0]>u�] 5=�����6n���u�,����\�F���3t�}�D�|{i�7�z_k�U '#���%`�|�y'�Ÿ]���d*�qarp4pQ��w\�l��6�p%�ؔ��K�coY���x��n$F��)��Y�o�o�t=[�8<3���tTX�����߄�)��ɨ]��&�y����e��e��U��DB1�"�����{�
�s�%ʨ�ͩl��K~�t�����|�i���9��S,qi��k[c�s�M���(�҃����Ձ@=o�L_��=�j?�?�tzM��>^^p�ƱLMT�:�G��\ЬT��Y�)መ��ȹ�;$�0�Y��cS�U�A����ev�|d�����~9�۸2ψ�<�1��_���p&����% W���C�CHh]m`R�
�lk{��c��P�I`Mԥ�b���''?3��	��e�W�/�
�P�B�b��w�\��(w��!b �5eĥ�m �~��;��d�f룡7��A�蘗]�S�Z6�O<�x�%�,{�m-?q�зi��+���{�,�5�T��%����o�e](*\�ҼןHO�Yd�i�=8���J�d~ �:�A��w�M�p�=�O�aՏ��y.\,�G�N�n�^��C� x���Ϯ7�����a�t�}ܹ�Xt�а%�U���S�j�2���z������Z_)a����gORpGUJ�_�
R��#zH�.�?\qp����F/*�H�m��#��av����ǎ ۏ�(q!Ǆ��u���,��ǁ��M�М[�؛(]}�Ӄ��T��&���H#�k�/�%K�o�r��/8*ZH���@ੲ5e�����f{���g��qlO�6�h�{��	&-�v�e] �6�!�`l�.r��G����N�GLr��]}��"�V�8����~|L�>��TYw�Qu�h��I'*�e-̫�F��ql��{�Vg栄��:T��m���;�:�����zG�/a걝����`�y�ή�~�E?�(�1lk�
�6B�����8Xhm�MF�Ȫ�>e��C��� O���λ���t�]H�5���S���ڑ�yn!� o"�J��J%��{�48��1T��c5�O�I���W�T�v�a�T'����r�3����;_g.�~b$�zݯ�L̸�� mb�y_����&4�<��qDS!m]R��q|XxA�)���Z�hޘ=�l���D{# lOC,T�GW��A@';̠�����+�7�@��*K���ў�E!�,�~�R~1�GW(����-g9��)[g[��&���~�k�|��v���mBb����-�vm�CQg� ��Lr��4��"��e{6�P	�g8B&���-�me��!?
ӳ�=�IZ�&F䈟};L���m��(���n��b��u]���Z�UQ;>JzmΉ��_D�D�ւ0y�o����HQV�4)Z���������:�P�¥7��lE�U��&-��#ڠPe���U쩄�� *,(��mo��;�����I���[�X��gA� g+��� ҝ�����k��H�Lmz��`�5�Iȉ��H6�Q��ռ�Pԍ����W~riXQeM�]�Zu*xV��Pz_�z�ak�xaа&�ւ镚�\ws�p�gu{�@G<�8(�10�)Y��qe,�������Đ�`�M�!ܫ��B]	4ĪP�8@Pk���%�w�w��4�I����t�+�>�7+�>���t|c�}��X�ϔ����eJ�!wA��kF;��5��W�?��;�(���VgZ��Q$ְ+ԍ���2��W�K�B�����U�VF�Bd�Z<��B�3��X��{� a���v���|o����U2>8��cA�c�V�C���Yc�;5j�����d�#[G�@)�n��)MM4ݕR��N�Q*���;�(X�y ~}�������a=č��#�6��5���%kW7�H��`�T��6��@�%�6���Uz̒� �_݇w��O��q3���LV�6R1�m�a�_�å9 �3�_0y���<B6�5�u%�N^>���!8��(�׉��Ԋ��	y�t��7c��G�&�ɲ���([=����l�,u�xe�q!��x�5w�o�eܷ�$eޫ1�"��V��e��1��X1�N�=�ɻ�B��ggr�n'ƺ�C�l���q�0���0�4��6j�H�bx{h�k����"�-K��J��!��{�|A�cI%k昦��5��`���Vs�Ƹ�T��/؛��3|a�����y�(��Ż�"N�]���̒1��`9T4\;p#���zp%>��rV�dV��C�����dr6���i&{X����@�,r%�a�ɾ�����V�x�4g�`��N(&�+u8�R��xS��.��=pB�ɢ���3�ci���� �w	Z^�"��8�ޙ��W��]`�Pd�c|O@R^����۩�:�y�-4�$ �>8��t7�[ZL�>>��3ơ)h*����G� 
q��S�+d����Ɍ�0o4��_bF&*���}����8�����9]�Tx2��r����ű9�X�*�G��iRG,R��9>{H���=�G����� ����%����|�g9c_�	:����*�}�d��Nw��F�J�fn���.�9l��40��j�UP�M��5�������&��mf]9\ZZQ�PJf��v�Y��_���wb�o)�Q�'z��	�������H5�+&��T��x���|�6�V:|���~ru�~0)��z�_���Bg��;�VjOt#Y�E�RIל��QS����(U�.*Y��{(5D��Ua��8ȹC�٧�#_��,�}�E.)4��(����!�T-�g���&/\��Tk��:�X�=���q��6�^wa�V$3:��4UV<�S�֐���(jP B�X��E���Hs���?t�ņ��R�j��l����2 �^�SF�5([K?7VH�A�W��:��L�	?���oӓ7�b��<v���n}��i�5�Z����c͊��b�W}'��}��X��6�̒}w	տ�a��