// (C) 2001-2013 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 13.0sp1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
lS26V3TSy3xzet8JTpxedfFpkGTBQEJYox2Z/omljwTjjfxXH9xhVuMR0wRbZlVthUe45i5SoAA9
hWOfd19CJZX68stUIKWviCkK21H0aOi1V3K5OqEJlYBe4rN6Ey/oGR9Ck0pVzHJ0Zn4Aoxg3GdtX
NcHqhf9feE5OWokw4C3h48nYmx9P1CTIkkmFRVtBcGrN2Bf8dfF3iIH4U69+bl6k/GlnAzcaXsVZ
rzkn5FRAuG5dkAYrJSBBYb/IOTcu+6Fi8PfwaQXjVPjBP0vNbN2JQmJHnDqRRwKs32UXIzWnTAvv
buqL+3IijoBWTiE6muzOTwf5wWf8B3qOK++BcA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
SGRQMU58bmkSF+XKMApbpezkdhGEpmJe4GyeMwjkIWopZ4Svy7701co7+lYsL5kswB8oSHD/xe3+
jACVUD//8/YL4BiDNY3MumkmPfuN6TfSAQakbpssuI1Er/hvPd+LvHItBiT9MHSDDLU/la9D1klH
1faRmyLA3qzz1FXRQ2JPPWvgloqiFm29jl1cJEIMRasunYFgLvv+wTTI+uE7pYhE9eyD1j4gE8tr
7qsLL3FdHkbjiA1KwK4MLt24NkOFcMeBJkZ5pot8GY5LTqjHkagHr1PTqJQTQ1fRtAaNIz7stnEY
capUUzjv/es5LyQPtmP8am6c+BNV5Lht/nDbEOZBuzmmP5Mrtf95KFeTBwgkqmtIh2t5tbj++db7
ZogOJKQA/2cItoVUTvupu1/7jrvwstTrD4VY5W7yb47AAJ3Wk7Ii42lHtx1BAm4r5jHb5Iwwqvko
GBN93boqcF5C+BiDd4+60+U4NLj1XACM+GI4VDyO0VE91DnjxTkLgmDEehbx4RGCb9e8ycaJs7WF
0uuuhsnmbV2yP9UUM3MeV+XdWmjjmuVSZ33Zsk98+cdJcLwMLWH+stZPP2albdHIQ5V9/gR+2GnB
NCN9SCNas6fYbXhlY3ydIxn18kx4zobTJqTn6luS88iqXWARNYT0vnxbjQbATugjYfb9kfDZCT08
J2OKCPgHHCw4+1BqTKZ5R6GGso3b2cW//1n8aJUj06iDh8cwP5Uwqbi8wF0Qm0mASI5hqC4Zvije
TTTlX78Re23pQoKY/rFUfaaATDvhKdNy0knlpgIQF7l0IWcx76jzduGKOtZWRY7kQjuJXDxZ6g/s
K47hXtr2SSwT8Sc6gKi4UYF+AiuogYW8fGVb7t/+omYAlDKl3oh98VOXHZbO02RbUZ8WchmLEH2e
Lum7qtqwzlTemYal0N4r0LwIcNpltlrQDvei7rkbE4NOjzDl1r7B0WRIUqAUnpqoHSzh6Szxrqyd
7wA6oVynGst/XoC6pWgbXZ3Y0db/cDpoN7jXX05EjZJWTvzrXoQle12+kWvMivhQxkU9QKtKWwQ1
BbY0/HW72oDG2yR6b6M2n/C9SvrP5Majy11TlXsZ8ABWkQd+uC9V94NIuAdGRDGr6tPWwseHJanI
TvnCz1a6ODPQ651+6giHjlpHlyZwlg661MRMYrLUt2z6v5Dm+UMkNMX54nDOM3NE3bmAUFPINQOn
pjvzEMfSl7UFNKvjXH0pVAJ57kmTrSWkfv8pjI6mj63Xt74j1LObcARpsQBTl/RsrrQqFQhOgvYW
DaX1eBlZ5YvRiZK9jkKWBIgZk0cbIAMKx8UlBK+Cm8F2V41ztJbqCtSQTAl7D+OxbUeyq+sU4T9M
dP6ClToBQocrWrDjANlA3FTKViiI/w0ZHZorTnFWLqX+oD1nQp+7MPfJyH5Ipy8xVjsWycL13olf
x/PR5zc7GfJgEt/+ZHojzIFs8Z5q6Y5jdUkSleMoqQ/iXPzBUD+maODHmKLPnYKBOdi2IMVjtLog
FdffgSBsvTREE/sfB/byTDKmLhUn2PEkFzNW+lFd5F5JO60sbqsHetchbB3J0DLdjkeyqRiq0JBX
CkZzA9Joe1NIIZ+sMc6rKdBUk3Pf9IOhrYd+Kn1sL+nTR4e/K13ZVcDc7QjCQvjukwDTQToV6/Si
UXTcrh6aXy10HRlGUH/p8nq53CvLF6n9VeZ6lA5K3YInafOsKJ3XScDM0vYMHxgzE5qtxIs8DIcg
/bJLYHbAZkv25B9OgSAArR9PyUyjKilqXFQNGVQ3PGJheV3c4CbrKx53dgF2hlm3PjETWAz8BR4+
dmurR8lo4rQD2XrEq/brEFIcbBwKMpoDAh0GL+ge3pMFy6w88T2vyp6iA94mLmPR1/NWKciyS6Ol
N8if8pDHXHAq6F9tWYgiZIzV5HHhLcY/PZ5GNrlubgjjpRD1FmWpcFWLspsDu216ToQaq6qKO4iQ
MB8srhta82SC3awivWSr2O839tSc2w6WYtbSAG3KQ3M0FmECFL3GyAloHVNDUhDs2UZ0TZx4/NJb
hYE0k68ILEcoLhrR3MBvYzHguekq3izTJwv2AvZLdOJd3owY7RkA3XK5jnDVWSO5RLfiVZEzhG3T
EQSkQ4QdSS/Cm5Yze+Uh91I7ZdlBN27s7vr+Rfn54jLGbQv3D16EEQgNPIqzUykTkAT1GUdZPlID
XNxt95C3Bs4E8ldr7Gnk/Ppjrh5g08iJiseoFubJl0r6NPTMQgLfx6ZndxCSjflI7XeIDxi4QDL0
YEJz8Pd+kaZrjrLjeTNtbaxLrJ6nqTMOY9Hv5TP0lMkiyyKiinCpb218hcBqq+BTjZQtecZFpzxC
d2D2TyZsEHNIhWiOXb6FTLDxbKCZeMT/dOfoKQI4KFNelQaxbFPbAnnFvL1/yAJtDqpVwoM4XJvc
48eo5zinUoi9D5IjSkTZe3Arp3q1448zpAMW3KQgxigbIk3E1nqSZQpXuI49sIzLeJmOUJ7J6lph
qpsxh7Hj7hxMx3InJcEgIMalWiPBOhW+sjQvf3Hq1zjRUwv+aqAhuRc9n4lKflyTW7acdj8HviPI
0CtmD5ZlI59Db2TdT1qhzc5WlSw37FlOT03V1RZzhEjlKbPDv+BtRb+gISukpJ5lG0S+0DRj4gi6
NzqKGU8BknEKX/6PNg5ozcru/3xsNk/WsNlwNGkIDgMhGTYYdN0+0R6Q/MzMWg91FuqDi9ANEJ4P
p+q1BMpV/S+Eh3h9cn3JQx9Lr2VEpotlhmXY5crTPzleft9Ro7xDYGJOBdFOVhUATKpEYy9PqqUy
NC/kvxTmy9z1AmGr9LGf/jDgSzJeC+x9QBqoJMeqmEyevHsqahafBFOnA6PA3AjrEeeQ95LizLR2
SLV2GLamE0H5k34jMKQQy2l8couK5DGnyLQP15VbICDwM4gcWRDx8A+htQOVzBcdNE1B2Ujx7peS
MV/zQVJ17BB1sr7G2nzPh4oWBtH29BMATpYP/WPvK1OW90g8U0dunZj+XzOBvXlDfQgjwzwSJMxc
hZZNYdTepgzuLEAzjwGxbIK0wI6U76kOrjpwNua/ikzHdnwA3MOYpuIbfK8yeBOhVmeVwMmzt6/c
XVJq51crtQ32SuQYEE4hHCYniHSo9C3l2oQhjP38n5YifaVqrdGUlq5fcB7jo+KoqRiEsa1bQh29
kD1l8JHy7+FF2Pq9leDYRzNTNFKO6cpZYhD7bFA3ElUE1jP6VNYpNAwKkFvoHJjQr97BrOC8uNlE
9lxMD+FpxobYyIbUzTJkFvC8Uf7popQLlfxgsEJJGHiR6BZ1vV4Kdx+VfI2eFaUH9eR//fHke3dv
rJ1ATQfijT+8oWdeY7SjDxcD6tI7fYq3Dvx4wNA4ytvlRrtaOh4CwS7B40MYwVwiudRll7hZwMk8
7hlauIb9I32jiRUc8KtPvDjzGhme0cMLGtzgGKhA6c42KMZ9YYxh4zW4YaH1W173jaFREWaki7+M
WF8nZQPyTuQvYfRi88SwrlZNlYEFimb5b9AYw6+PawRi1haC8eAhEPlnw/Xt/FVIbKnA0z/KdcDh
IV2s/2h8cfRzYo7nAy1HIVPg6I0I2uEX1flhJozBBqxCoANh5bkpZam0yg0utQwJ6OwmfdNSTOW8
kyuKPzdVKJ39F4MYjQHMpRL6OpSP1IoGhn2R0Dz+HTH/qK7rXq0AF7b9vT2jRySxs35RBRzul5zE
V40//1OFK2LQg5lcx+HkydUdutklLNnvxF6k4Vz8JH46G0CSh5TMMaARkP6nViYQ8K5uB6it1xW6
2JKh0Svcyme7F5COvBT9jtijFUAJgo5l5Tkk5lSwm9qMuKN4/cnAfBONRpdvPjHc9C9TNUKPXRU9
fhPu2OP8r7ljutOc3Z21YNP8tP0Ui3UsfziPB3up+7l2eSGUjgolYkUA5RBtTef+y9rs+3vVjhIM
EM+NkQ9ltH1gqmBQkV0CiQ4R7XdxNWnHhcQqqHZQIHAgLG5dxsLr43kkx+/Wp4uYJvDhLVC1VAcD
2540qixlmcwYVAbW33lX/6ooYpQmbGIsvC5tdEidpQ/WdHqkno30tWWH0Ov40KX3uVXN5WfLmTST
d/1TrztDshauMz4JI4pRau6JT+yaK/95SHHrqJJ1lmIKz1ZkM/NO9sJl9PPKrLLwCq+1AxiSi757
0P6Sl9sPO41YOd9JK/2zlvR8top1asfuJOhwNwLKck4tMxLEd7Xd+0TcE/4NiX8DyCc9f4M7DV4h
RH2UmqgzFjDHHgJxtuWcWJCQlKAFvbU7vhAbQ0BSDy7IskG0/cRSQzA3TLGlNNVdfVRu5tKNyy6o
HtC6KAwScwBKtNNeFXz/X7VFK9SLjwvok57fAMcb65hmyuA/gmXt19BTF4bfe51Nfy6VUoO8EW+h
wFnJZvaacOCPSoF2luGFFMr4bfV/9eVh5xkTBcpJgqVGdECHygqOXx3leZYRrLCoDU4zBFhswAw8
aTfyzmFCEztTbcfu6EicuYzxzMLmgRBq64qqZzUV39FWSDt8FUdmiDheHUVEfbK8E7+XIKD2o6nj
9Yrn69RFgoB7w8zef8p51ePVwu1CI3seP3uZfS8hj4/05OVVQurm6E++7LJJDCUeKHsV7LpQm2tC
7aPEOeF69hRZ5KaP9hYRTm4L19MFWjxXp4L2Xmhop7qGOXbElOBjsfjnCV5gdyuNFJkTsj4tDgX0
ZnI8OpzAm9zkvTVCFLH6FS4lAakLv86qsK+iQMHWHYmJmCJVYB7jB/7NJ7uVq7+cLwUYHIT15ZMz
EqylLcCWzUhauykphf9w7LNUKvbemzZ0pJd91RN89wsEPexpYWUeTZDif9+8+6upg5xyK3wU+Zic
VKDUIieQuLD6n2DOQSJkIhVHkw5yMdS9ErZ5h5v8mS18VRXxWBKS2YXYGeTlwvTVZifQUvP/G7PE
gLVVfP1PrFVWHjnEi42zl2FhpKuhUpnWkmqZugI+075rNE4+B6xn0OPBYKGEIzqLMa9M2h7ACcyx
d9hF81ziDR3SbwKtHBtcFSk20nf4fcAg3HB3tGflyTH6zoqMIb8WOamhDbCRSV0xQ5Ghmserg9p2
6pASj+bVT68JIXCAGljJ0GsNkNcSp9aBHOC0R7L9HvP7sYjzCfWCMSqjnpdJsF0eQEqSZFwXvFJP
URej0qQOvhA2hayl5WDccBKwLtFVI6yFjYGDTEDS8zO1bJjo4DdfhX5CGYPVdARnZGokWVPlyWzi
ybzrqajVGLGSzXbGAu4eU6LwHvdMYODkE8V5FZRZuGLCd9EQH3xIAibfbjNT9R7OBkSZwuRZImIP
6EpljTrmZ4q6cTwvTUsa/S+xekv5fw6USbA127ID3bpshwFJSY92I6U/xZJiVBg5d9Mb87gm+euF
WUtDWzVBtMH06WGGpWq0Ql+4+ToStFFRI8VGu70lYm2890s22izP+sYEunOUTmDehlxYKkg9QBYz
ZpZd6QGFlpQuZeW4E6zttsaOL0jhsroPL4a+6tUltnaPlZSENoO8MsnPu0W+MlSyKExpKw2XR9Ci
WbJL1HrxL4p26jSj2adOsPIjA3GaC81rdlc4RH0pRAP9ox5QxO7Sd0pFxT3IQ8Z22vtPkspfuSB/
dBvhNcyG+M4ujy+o43zBhx8XDZ4fpaHb9RG2NlpUZFcI48O/A9O+3cXbkmFFMOnpsnnks7Qh5T3X
k3dcYhXDdRkPkoIEqasxix771Ycl9pzS9L1+rCHnLv9mQSvl9jeNMDqCbnuRTJJ99lHkTQJdQhbW
RV8T20sFxxKOAHBZelK4646x17+ARwhJFkQ3MKRbnRFN6lNbMzCa709ntA4ehBIrBsd7N3MYJ8gf
jdj+fUeBu/LUFEb2JK4IOLF8o60BtnakwJspGu5h8hjag/fcMFztuC49qtsMuO1nysryP1VJ2Aub
nWu67KozY5K9wkfq/zauxsjW2KpVC/LoE1Wvi1W5XKAM/7sawRJ7cY1xdL0lLYzMM6qnCgaXkKjm
8/Elt3F1tKWvsCapwrDIKo1IJfvTcuWeTFSRWsok5l5C+QlwoQ0e5bk0/mAYB9WsBauE2VJ+mA5w
MegKBU0Kd2Bud0tds9xTIVBC9iVJGB8ScfEXNxil2ruVY+jnhhf/UgVbWT6RFpNjX8FMSSGouV0D
ga83MOC9XIHeSGWQ3Pl+bZa+uWAos+6ex69ymP1RCR5+loM5wCVPLjuKwbAzUcnvhB9Da/8l/P1k
ASGHODORzWj0nryQ8TyrR3GOzy9lSPSZeUPUZ86o1zITDUPX0gNQCLmtrHqPvdGTAWWjYu7R4iuj
pJdYMEOIVe9ckKgPiiHGnj2bwh39sRhvk3CYgJ1fEA3Tyq+o8ftzdENQFLK0m1/SVrg2xM6l/6Yh
G7vyxFNVJySmnOEc/azUoWiyhYSwQB2IgVYcU4PN/Q3VTHuM11xC5OLKX/IsvwoXPe5StobqjRJV
jXaYHgBAZzQsvCIXTKtmxboZ73J6vxNemo0Hby1nrlcGpztN3br301xMLPQuN7CVx0FBW4uCGhPI
Hxa5vUUYxID9ZJrltxi2oDdNKsWuvZHg/j3jToLu/2fs3jRXoVuFf27zG9hPNgPZo40bxyjavcMh
oQc/42wESfH47UKmlKNkt/CeYkyqxs4A9CPhdT0IHvtLL9fCyPRr/CjAAcAOQg+8/gQbh4634P2S
zdDPYs8AZRV/lYP/DNsqVWTndR/Kv7Sjc8z0MbLBURfGNeY5vcjELMwAC/rdhPRkvl3d8sgWkn1u
+7bixoMuHUh6uY7n9y1YPY9+PG8Mg03/EwLnBZCGJ3Bs3VeB2AaX8I4Wh7SVnqGb2yCzN/Xt/Rwj
j15jmNFRgnYMuFhZtNpeWWVi1OWH6yd3BzHcurhNEEF3Es3xaZWKdEhFwfKZEh8f0LhY3LJ/nhhM
PSo4bSvwq9ZkftbUpufJzDcwQ1VIUXVve6Ghm/XadPHSlNksH4KE2WxowN95G13MFnJfW50+sUaS
srR4uMK3oAlFSMmWz/6LutTBBjLwhpTQyRdRQdT/YJ4RxoaUOgr3INT8ha8+Qt//nxAD4qN9lGDP
VNZmzetpHowpZOkIFh1WAhCd2dgpPsYpeemJ8cKEwfeV/03ul7XBUwbDkVcoK50gAqnqt2e4BLic
sTCKU8H7/CPzrQukchXMy8k8nEABn/XNCBMAWOIWm3i45D4sxB0JZvyuIL4xcRTpwXgnQdGb0Glt
4rsqq/VtpEaZWRGObQQHJAPCaPRH72OXkU+vgMkM5GDQK4r1Kth7ERZ8VOJJJk7eMiDslX/OP2DU
zFSEqCOIqFzvWDK7Gefy3HmnnadF3zW80wVGBinO48bAnV1cpWwbYshsylWPXPrYt1gSjRucA9ry
AcxpV58qTmo7PQjLen16PJS1t6Dl2lh2HCgnWHYZtFlPoJw7/qCbf7EyAbGmVR8n8Zy6hIPyDY4s
ioiJWMeDKfpQLhizpYphbvlmreJzAVK7BpN6KqjEo+v7TzG1YHMLg3vZ1JbPySE0sleQpr/Opxx3
QwgDS9O7fagg6w1uJ/Hc+F4VR/zBtbJuALO9glZfUe9u40EWjSIgIQJZ0vi2U6IiEOFNUywGIcND
IIxOMrxPjaF84BjJl/peCBzE3lctrS9Taks6/L3YQ2+wo+A9UY+v0K7PjRjEd5YQUHaTVIS9I4ky
zMEkOTn3ggS4CMv4Bn1CCxUSje+id9zu6LmOXf9e3vlOljr7oL6hrGJf2i/Q+7kUKzxeIICMHJrq
L/I3wF4c6bBXcIsQcxhGizEdYyN5fT7mhWFthjJl5TD5/N7kBikqU5FXmq4SgE51UmoAQrsPAxtj
nSIYS8hH6OVXLN8hpwRaa4PZ/JhpLR90+CYGhrghJu+N/jZRIpIGbU9NgwAXuQJ5mxnJrAlRnVWb
+JYEO9c5Tok8fXglQc/oLhkQT7mYhhCYLQnXULHD1fT8QoaODC5dpFRVsXEF9fmissgRSsEUqyXW
nSWqtVNcW6sQnFUssk81OZtf8BzJrIJGj5NJDsChLKoFq1e6s2wEGSGy90t2Nz9QLeFB3uaUfPbZ
outjGoL7G/YEO18T7rZQWDX0HiTyPhA4yWNXvCsgoXMX8Jqugu5d0Wqfuo1mckmrlMHpqxM5hPG+
56gecW2YltkFlOaHqZ9+Dw/Lx9Z8wnElVDVt1k+qFZMYxhG2Q6BdQ6PRFAUlQDhR9vxdRMAduHaC
qy9lp0NxVj96o5+BSCVuVkQ23n7ho2nRu2YBafXy3I1ax+erGKQ0Toaym8Twc9gfZOvuFVqobrsa
/xfgNeOTxHGk0mdNG7JKoq9LobUwRu5EpUyEBSQGxNzD2pEXv2tfMRtLprhrS3yoXzhNCD0jLDy+
NB0/sBlcq2jmGTKHP+P0etsznmWoJbm/2ojgxQeclIdgmayhngmA4XP1kzoGLHM04ZKbYboPe4JL
TevG9inIClnSZCJozZU2raVhONaYEqVuH67w4uCiYBKW49TkDiinsFR/XrCRIb4R8UVtgQi6uw7F
EcRGOzJi2HPzR15PQ4wls0fsmOQ5QGiqFFRvxKvm9lrbB92JhEx7oIFtSfGJCJ5O2w6q7Bna7WJG
G/Iy6rFjNZJx0lsSTDC3CQt/A5ZqECsToLAwzfu2VENYTR7Xmo7MOZLMaGP3FwyRXzki/vg4o3AQ
BORfb+vRbyJyny0t/Lzihm7Yt5/VX9HgSPtmeyVHmnX/SxKA3Kbn32hb/9DgiiNZLGtXgrUi/Yi1
TKRQYLaJfA9AnnZeVGj4qey3gSglIQAqYKc6FZ6I+h8kcQyGElMUdXq6nnFrMTIcXNtqEVZ2RKL9
6BZQX+gBKxo/gYW5fqfAxN6zjP8QtRZTSpUiVm0/3VkDsKUUzSdaLqNxj9wrOwyMuiia5Q1XirSP
7HS77guX1tT7HPsUb502OASBfnkfVeYP5kAevsX4hqihDFGHleXlksulP77Nvq9F8m5GmZnD6gzN
xahCIbXjEPGZWyuTHdLVXJueR384g9lOiirBs+uIMTl+69QQ0e6Xg5G45EBCrx+vNwJS3bUI2Mqb
df97Dbg+FUheCfihcPhKOv01NJrSPwHvWcvUKu+/Vj+uMT3MRq2aGpo/oQUTC0BmibFqlW1pvzr1
XY7Xueoz/j1eDBhk9GA20L5eBy66ea2vIwyn4ONqnkluF40Ngw6B4Ifxspi6mUlNkzpYaq3g4kCx
QjMmhFJLenBm5PJ0SoXwp9uRSS2h674H5bNXAbUEY+F51UG0nZOB+u6OcUXxOB6NVdDk4OUUoZOf
Dabz9rZfWTDeuXtjYFBPo6fjJAD8zL/HMc9L4ZgvutVWwcc9qkbQ0pw7OUILYEeQPP1eX0YvBx1F
duWG1J8OcOIQaDLZKT0D81w46LOvlzQuoUhNIHaTTVDviyh19dhEJaE5wh7+OfHFlRxOagS7HRUT
CaYKabGUdLZtQ+zVDtgmvH4g91ZJ1FmZ/jxFjbNPyFxST6YBLBepBzcCjv10TeBw9pC1tUAyavsV
+CETvIJJ0zJJWSbpfNOIg/Uf1rpowO+AGP9+LsnogA585mtqdF2kll7a1YOTLWI61FBLgZGnw/84
CMhUcBUj/pF3cBAhHD7CVCXbO/IWBpHLV8GWyhnQgLwX5zeGDKVHHECsPqvStmGGl8G1yNLfjWjW
OzQb7QUdpsW1ORlw7MEE0FJWy6Cbc1mvyOJoiLTjAQ511NddC+akaC+40DNcubYmTu1NG8reQYo1
OLcRpkSV++VwCW6S61T5/6oUv4XG5HfHHDxss58cBCalMqYvAXfTF4vfFXxxwEeQHE2pDjz0zmLJ
iqCXpN/Nxj+LOLjx/ydX7ZmnfQy8fA+eKCPP97pNCAV8Ek6lK2XxF69z+t9pNqk2Y1nQCudEzOL8
yaCB/1w6A9RIQXFHGR2N8NSEuvFrL+vLO4Pb/kJ1/evDLobtotIvti9Zta7uwk7zkZtP5jJ6BC3a
UIxLRzOMlUfWsUr6RXl66rCJz55A6YuNIcggbbp0t+VGaNgHzn5j3IBbHqeh0Rb3Sm5cgLrRJ28Y
ih8+pfgMqhFt5nINQtWj6Du0LSmwpIQ/Qp43IHPZq7XCCWXbs65LZrUMadvXYfdmhqGHx2UZhHpV
tkNjZelk8xHl2HObyCCtBpN9H+YbV2lUu9DYT37KrEROcyThcAPnBDaEep+TAiiW/oNW0/xnKpGp
0ioNV1BxUqD4S48Pp6NP1Kzm9yI6/pNRc/GFgWZx0Udpf9giGbvJ1o+q7zjLIueoqBeaEM2Zs8ko
6LjLYqGWdXDtg4TmJOnTr75MgUweuF8aKGRt/oEQKGI3dWU/Spsl+QBcJQEP/osXDLCGaK01d80c
wRs/Z5eQGvO/PEQnWe6t7WnDoRuWhPHEo7KmWYGKOKzmGgXrhhWRjd1gVu4EXuIM6b0L1ggw2S6B
3pQ1GhJmLHczpn3EsZL3nW7WTH12IXw9I2gYe6EKAlSyNknNfMVj9h102+d4VjTmM9k/DW3aRkVS
zIFwYj2M8l/icXw10+WjaXM2lGX2BAeSqAgGUGrYhRa4NOjBAPIRvmDMdpAHC5oZn3xv422UrmAz
TYKhTabLPbK5Hx95gFucwVuDeBVUTWh6uNODMW6vMClrJy7G8FkSuZeHyYgP+AxEHmlxnlua90Qx
80QMQ2yofhpHNgjhsA0WgRjSB0L3S8074rZyC8obzyWSCXZEgS3KaxX7mTiO/w30eaGQk1v1NOmn
7O5oDX3RJtqwhkdQ9dLQgu/8sYs9Ts5c4XdaDwjLqgK/1lpHE956iWOrXw9136JU41xPAoBgcRoE
NF/lw+u6jF7x6KzlotGKgyxZDi9DLRWD4UDUw3Tulh//9OH8uBUjB86rNzAr4if25TQ7U8kvqgN2
b/s7BAnfQy4ec/a3uYDb3qmDVCzZy6VkaO0nqP4RJzvRtFjNNYf7MzkkoZPoJbYB9Vhmjvse0XR/
W+6lvjYvIb4HwtUP5fNSUc1HSn2+1oMaJE3I5gkjfPVOhOrm8Xx1klQeaW9Efl/eB8wApAJjebod
o47j6U+jMFhzsgyC+Dl4uzXRN5JYN4OHYs53qRDGPIFepB+IlztGoTqHMMmOdgchKWctbfmOiZAS
Gy4vDnefiGMY4Ys9+nCwJT4JbyJkTjYs2GqEekhIjBMP8tPeZ8iUddJeWRnonRkZoBmx68Ec+fjx
2U0gINvX/yjqseLNIfc4bvAreE9KzjR81muRE/CrS6fGoPHwFez9kzPFblsCcdCfqliAJ0wg17D+
4hEUxqf+U3BQXOYZZeKGh5nDANwZ9yNO+YmKU+5ElwTLnWr+CW82azx9KMdE9E5NjIDAQte3VC1f
MoJZM6q6MM9jeGOWXddzSuSz9EgQMzpVvBLsKgQWVr4sLSLfAFhk+NwFr/e7SgEpRaplXpw+Y+fo
TaqW51dFGKjOdSxCi2TDhVnZmGSQa7oFCVwHtaBPRHbITU+sYDhrwE4wUbCL0cBMlFfaFAkFP/ju
WU2CtTSxCiG5PYkK3yunzTjuCSTaKsiD/im3+bg9WB+N3oepe8MEBwSNfY8k9zt5i9ls0D5Jgy4q
ulglwbxXaEo7u86L0VxTsYEgrOhhWcqtzK9zlf+Xl8z8vTajYbZdtNeBIEoaa9zFudQUEPmZcJTY
A+F6FUicRj97Qxpr+g3Dnq2rV1cOFDHApUlgNiKkOSo0+R9XwZapJnB/S1nyES6zHksK6Ii0fZ2z
dci7jdjQxqk4HM74aBtv/lZx8roG9r0hvmmNOMn6FyH45eVN2UUJCVeOZXq1IG6g5ln+sWSLPB2Y
aQMcp6BbXSeHKIEGkvWQhl3gQrwJeLLP313AER5WzQZ13QO68TFgLyMhgK5gyM+9lsdQw75UOjUk
9sWnRJLuAMhl4cn0hwe4GRx2bFSqEXvhPOxL+ZiJqVrKhjsWpQJId3VzfkczpFa5agc9yH3R4wfe
jdX4J4+n2yHsJ09QhqgZ//whPMLtA0a8qxKzgDtecREimOUirHtZtGF3a7ZkAnyrEKCMc3unprAE
ppxw7U24y2UOI7iQIMCRpFHcC7z6nIbsZC84csKUjDl+HB/r3bu+XvCpzBrI2i4G9DCDTTboPfVu
4EFaNLegVCn0dkqlzSbsYYZUyoBZqB0lpAXaFNzSrFZXnvrxC+6GgR4WEgbZU6EcoTJRrO/R35Tc
B94g0+Yc2710JmtF6RsCvt74ogFsGWjst0JuCUMK/bhuvlN9pPhGN9uOQq7hDWQbAcZIWH1g9sKl
he2Ow2OvjAaJ6ibkgqCLTLcBExnVKOIKV2AnxxdOsRbtuPRphq7Qwf6axLKe5Ticu7fv73Mzoi3Y
vTHygxmV1zHwKgptZbzh17vg1ibQAWUj1DEYk7bja1G/rRgdo4aDz/eMq1PL2XPZfXocVfbvhXLA
r+ZEx8tW7pdFjgIqGtQWEtjA43yapwUnmDdG3qyUQg72yf2H1EeaOJN9xUmMPjkXMc/N+G0IBC2I
lOepQetxzCNqY9AwPl3/qb/mvPGWYHNvO5rPssBNFnzLIz/WHbOVFnYu4Uq8jgfDFA8p9Bn8ATCm
QQSsrPo8+Kn1iONp5VcEg9/6GfLgWvSfCnVvYQOlKLEiSjZUjpLHPqtWWTaTeR8zPJae5kSl2f9+
YmN+hCQ25d/Hp4i6wakabdGWhWDYOOZMilfe4d6R1x/U7h2Pk0oocmjATWVXMiSHk49J/0CLM2vh
rFKE9Nz/tf/r8eQwhOhG6JFzAJXb9VE+CWhx40FA9bDJz/R52DtxqbLb9pPTUegDJYiBMU9LQwKx
fQ45Hdxq/5WGkiNJN7J4b6eXO+51jAz5hloAkdJdUoYVI5oAms5SrV0iEvYb4+hVr0x7PpNi1+Ka
FfG4T057VpOFLtQhSGY7KlWZz4yellL8SEv4F4wza+PxwiEiv8SJt3YhC/9zbiHeOjbYFD5FoAXt
osgf8gsiKgg1dP7WBM4tS0HmNJjkresYDh1R9V6kmlgIrwHJybwm1HgTZvyg2P9WIfTQe7+Dl4Rq
Fn7ds8FJJk8x6XcoqLyvdLDtUhm/JQv7mZjFXwm6TbEW/EsOpvaCwZhPT85xzsAEGnRcHX30/f6e
stbE3AzuFFKxGrsZsCIL9a1b1w22acaZlk2Gow7deaoKgVYJXi+Q+7KIiezJJMIfZ0axcMj33Kxs
EQCTohcR8alID5HYCrsrlIzh0yE241+CRbvhRQeE5JopVAoqJi+z59/SQU04RBG1RW3P/pk0fNPP
oexD/JVt74KDqpqqmp6VNm7Rnmsd7FZusEGcWVTFUiV3Hs2JkvOsUCqUVVkt9LO9NCDFaw6jMfl4
vcqS8pmyS0Gq1xN4CPFYa2msFfbbEeeI5gFAIy5p0OgdV+JrlEVrk7gjbG4JYqcjJoVq4mwTGWf6
EgA1QfL6Hm95/b381zBWg1XOWGLciztBAInUPKI35tQIguXnC0ZAOiLY6b/7uEef2BBrb13t1Bk7
rakN+w+Bz8t+WRy4lhR/H9Brq9si7h0za9KB8HqyHRoZxOYxDxVTYCGTezZ3rg+loH43kz1mVb4L
dHfGomMW2g/pIfRJ9E3plXZYFI2hBsWu8eBQLyVqSPcn67EouO+vQl3JrjDdM2122K6qIrvZ3Z0d
Vlo9hY+Nqg1umZnq7/3EnXVebRoA3oePu+Pk/ITG2vwqoG6iKE82hd5fRk9Lo291CM23+MEaYMaJ
emlrhcltP3Q+OR5u22zonDBrPWaI62Rrg0x7NJxLKuNmn7EGcg1NKCQa0OqBW/Zr/CvYSYFJx8Fm
rJSX8iMMQo9OrwOcupqtf0tQGFsXn2zCbAEx6sNuTrCqRO5/aFTb6dfMRsGS3A+g6jFB2Ipv4Si6
plGPXxEaNQCTO2chDRO1IYAwgoTN2WXFJp4vdNE0PR8giylhn07RGhKlRQiLWTGMnW7ZvHRQzrNm
+GKMjGxyA4l0IInulqzciuBUOlCTiraJTQq+T4AUSUWcsv0CEiqkWM8yAIX3U9vl9tfA4lQRHTkB
uGSBkfZEhcmiKLOv56Y0QXNZbkt+WjTNZ9unAklGWpKhieym5qGIcIFtYUy5pLWQ7A347elGIq2u
9U4ETUjhnlcv7TGQdk9yxOluxXqZnAB6HQKo/ZdAZ1GjKCzJWT4QkOl3rrFV1WvFMNbwGWXSIk6S
gA3Gvk5AI+9Sr9/FESRZ5rjgTrZTKC4jzB86D6Pdd09hZugZ0H+YX1P/u9XPz50E7S0cqyvV2zQz
w/dbtYPNtHhXqcDq32Vda9HlYkyo25k+9IdVQClDI+Iylp7RZZg8O28XwM0QtQIEaaCpGbijgFRN
NQSZvt+Zr8cUiT1MLTT3JHnR6X55mYuFC4amzikHGKhGLYXarNQLwWcnf5wHlvKcZMkxJdoJ+eCo
q3RU9V+B9A8sKF9k+FRQm09B+u7/JQYcxxcJa4u+wVP4hhVPWLtF8JBtNVX/WJ3+PugOA7n1chOh
GKruvIcUrS8GARy/RtPTYLS37rKPY7Vs5K2E3h57JAUVkhKuNkCtpPD0c/59GpAgw8gMeXtZvIMx
H85Ytm11si0sQQZJOamLd/BgD+ztxhH4E82ho3QPY8pt1HcHxvVnXZTWOQ51eFjOEbUKoev6SBKJ
2zPOU9GU4oImz5xdVETNEJYVLkPNNuVW+mDxIpeIP1ZJqb/aRSLCvLlQpPn0jeNa8MWRDOZ7d+xd
P+UUgMGtv+dHbqHlGaoe3pE9iy8n3/CJOra1trGn2LbUEWgINCOAtPScKErNs15gdl1OF3xZ12QZ
07D7Qb2+gaWJ24/h70qy+CoSDaEqPz+QOJsHd5022jqmha9F5+jrd2KnKFUQEhDw4+D4hbU7YeKF
QqyvrxOCSnOqHT/a+nmjB5czIScFAuHSznoxu2NSvngmY1MHQ9XspeTV5/eMvjfJXHqwYoznAIwD
69SAkheywnYN+2hsuhBgqdkISrO4K0ZX6OizOHl8PKQWJeir3nVroQoqUdD7buONkUuY6yqs73Xn
6pNFkrMmGKAS4aILGWTHGzqCEsF1Y4WclMTbAJl+B+uodeIpBwb5H7THKAZg3iJMDFqb8LA29JzQ
Fkjlm91rlBG2GRaX2OJYhUvWj/PuHhi946gyFC9I0LMAqKgTibIDtN1HXRWKKzHCoXRMX022SXlS
PI9LbvfLp2UWx2TK23YttQerFNJZGB9xNQ25cYT3IBWrlaKaVpdVnB2faICPBZjUZJFZ3OYP2jIZ
SvgdkeYoE79F2lDfIM7Lhl5Cjmvx1C1DLY+Sc7RwZL3/Z42csXoniswAh3ae2M+HQFMRvo+Y0QdF
pVlxhCUGKBzWyyCwFNK9GW1jPZzoQlITDBNvGEqayHccndQb1GZ28sIE2UfkKz1lGdkFvtI5Rgrc
jhUZywlJTABxDo2VB6LREKDoJes/pMAb+pvEbiYSGJmls2+3bSvc/5qRXrzSkNXeiX07ZGReNPih
Q2US2FjpyOKuo1K2AtccUVQewyQc09vB8x/JaqSx22H/bN/XAfiV27eCfau+8umrAgxJ1AABZUDE
qfTazfyJMnvGwZfa0O9yLMhTw5iGey4tmMMcXq1qRBwJBt4QqxlV/4nWzoH8hLd3JS1S4ES+YuoT
4SAdddLU6OdXERXkNm8xLNHVaSzVy5ufv+sTWCGI8t2SJSWvCiuJEaV3Wm0Pp8Bv9+q+CCgEvGUe
P+wmxSRMg4LMD3EjD1ZYQQioMD+gE9A7IMJ754R+3pNVWrCu5jHywtwjBvEwbcPy6mRTATGp/fBV
U1uPd/3HwPsvn7UCAnd75LF4eKzH/kQ0I4cs1zmPSVqhACTKRR10NoTPZ509Lmym1KyZDQJKR4Cp
xtEDnE3r1T6WKiZwedVX0vr91QoI+zvJAot4CEi/EBQe47hqbuq0c/w/bDI10AqE75K7KOSl5HO3
lDsJagahF2JL1cSDV7hIiDZSV/8anasWNI/ror546hmZe+rMDpAkjXprMHkd5rWa7K7MGeeFxto1
U8DS6v0gd0sjulI86rZbifc3eOt/Qz61q314b3psLJ/1bX6yUAipHhPOQ2cIOt+HOkg1Wu72vbVC
Ofh7e0SSSgT3dMRVPJTZKcm6Ho+JM6yT8QYVyEaHlI/4zHnczoLch+0+gb82bevs1LXtgVmDmcml
XkuPEqfqLXcmEsWflQQngF9pRpKk8Fo9b9e0JCiLMAFHlS0ir5bEHnWFSaC0cU7U4OH5BDdviOfL
OnNCYSaF0x4oJ5eYOfXrgnev6VYtKqz/eUKmNJklqo051Y0e/ablRgcgRvTC3nSc2MTbAK1Qs6Dx
2QjN3w+rBw5PKxKAj4GnYA866fPUSQyYJRRCINNXp7g6Npxw6RUw64wdD39EBCVxiz+LMQB5ZLcn
u4wMXr6QywGWuIG6phcNg7ndnWhZecikLcivVbfebVOySHoG0F5VY0UYIE5NhsH24DKbjYN2rfg3
7AcsUuDupXL3pT5d5HIq9gfGThfsoBe0MyvYeAm6sLYmpWKoxIAlj1d9qFg+w/i/VEw2PhsONZwf
W69wPpMj0RfXKNz/624ZpdhcaVCca57fUOOtx5rvYyS0CplVfbOyaGIXnmCEPZEeh/9s9V7RVvVC
udXi+XoBO7rLDrLtr4ZupbviaGn0E/NmZzgH112U5CPdmO7fDG8qfht9KtyVx5eoHqCtWy1+7ZTz
ST1nMjG9nhjCBBFycMEdn6C8OVvUKQUNZuilMSn4NSaFLT+J/IcpYalPWi3P8iQXMzGqHhmdeJSz
lVG9SyjVewkUHIyCRTcFHmo+eWAM7g807LDzXANaRiuGPvPPQMt2H7tRJDRdCudAC97ekoiC7i+p
J9UqFR2B3ffcOsGdJpC77ZwSHCorRl0wRnyz3GNqKHkyIJHHLsi0Zg3ieCoL7AcuPpM0Kttlpe1M
FTXdYJeztPhy2F273j8MtmPus3oLKvJyluodtSWosdkPb5rKkdkX1XSwVp0+kcEgXWe4F3SMDj4T
BjhASwLk+6SORo73C6W1M4BIy4okAFfgesflrlrqttIVpUrzbu1nROH268rZgUCXTL5zijxwKT6Z
JSHdoXP3hq5I4ebGgRBT5RuX3UbEVtQn0kcZMgW99XkeFVjqr3+62qBKC+dUwKP8+6C5Eke517P8
qVOBqVwZlBT5MZynGRbuVNfcVXVagZN6JRyu1A6n1uV3i9mCHuBmefG/E+fihIVSiSyAaWr9Weow
8lsW7WTensBexhcvcX7WmigWKDFcD6PmnMnZ8eqV0nHcwzjHvEZFqxl1I4FQclERm8Afq80sWGAT
JwGZLr/XUKdCUORNHB+aSN7U4DWJqGorMq0VQrVZMAEbk5l4EhT9TmUfUAJtD9EMZZnJMwxr6o3/
tU+PX9q/k+mcmA+ZGKHvwZsnW2Aotjl95ADI41o4wo+mOv63AFshXghLH5IJZoKYUeFl77VJIoiJ
nUUVdnB8TxeX4tmmIsFNksdaXVOEwb/ofhdylz/GTsIchqDEnHzQRw5GowO2bt9t7z8CY2EYfsVi
jYWnwa1Qyf3Ra5IBAvgVVdoO4cIeG6alTkEtTialbt6FTbUk8nYmS6RkirLKvfQjMsZUUYG/dmBn
W8nOR0vdf28MQgHGbMrcjVdAgLC2B9h5YMaxq3sfR+DrdO0jqLPU/r9PX7xiFPPa2FhnT4Xz1/Xe
LlogXKfhmj93jZvvh3Y/3ffWZU7KtZpCxxKBL0dWu3lC8yqgfR0mvuKwhflaZp9IXCeayTGG2vjU
5CyfrVX8ujLJyrR7u3br9bMx6avcHYJGaCpiaTKcHKQj51yxfTd5uXvoL8+Zggxxyj+jVFJ6zYiH
K2p+W2BXSGfh6Oxd/4rqm4Uv/wuDlvd1BEtck6kxpTZTTpF6oUjIBiNRsTnlM/QwZpzN/MpoRW65
K4C71bXXhUWvv5UHQKzA/5gizaUUl50RRq897IVbAnaFNXieHcyYE7zwksMRvqrSyXeVxhTWzJ7H
bGLf+d30JLY6RHKIbyoLdj5xmQGCMDLhN6gh7vDMxun7RHWRPvwKR1reCF5LSYsDIs7m8gor4/QW
gJAeyDLqbiXSHS/yN2rL1YRMGPPokFmPKmweyZ33+D+MEI9MLa5Iwuf160DAkzQPyWbdtF1hSPhT
beVVs8cOsUCBmkl224SXwiOqJPQx5zgJwVgPB7ZEeFDy1jcRozra319ZMHDf6RYwyeIeXO3+exPS
v8HnrMcL5bjLtrTcY4Jcg61uP3K+Wss/3YlD0NbneuT86lPTo1lICPsALhS+IPEhTDvbNJuEXuaK
W1AKkm0G440qasEi7JFh0dp+dnO/fbN4NzYvFMlvvNzpjZ72cT6N7TVdIGrWlao5UPip88jBQZ3Y
A9SBxHa5iEC5NPp7F+uKMPZO8VmIkDhpKn4ywXc9Gm2P6fdW712czBagyLidJ4mF4m902DeDUCP0
kqdR6enHVGA/oT9S2w13ywWAkSSg32whg4NJ6cUbLQBVl0oID+MEvUmSS3B38gbXO/PuxxJOcDwd
E75SghDV/bJrUKB0OSH7Gyt3ZTzjpPk/9CBJUjKCuIt/YdVZ04XeIW73mfhnsSZUIcrBhM2nOAVZ
VMidNeWpzMY9X7EB89zKwlEkGqE592jfrOMUVB7+x0nAUwjYjOe2C9PqWbRDWpmOoE3RiIY5wd8e
nMj26ukXvICwLyD2/hAJre537+T06niLe9F1xVtcGiHwrfgK01lL+mwzR3lMIUoCG3Ilhuhugs9v
MynoliOERbhx4Hhi4UBSi1ysrM2Lxn75PTtXaCC1UiwVmwyU427NlgJu4K4nNlKkt9R3tB3OioDv
fdcHp4pdK0BvRb8PfZf22qgXygnfEuKjePrhFImFlCcoI0kmJ8DYZ9j0UTRhTpEfFOH2Q7m8u01D
cnTZ/mJMmXGBUUyO/qihWSeRG8+JQNQnOXJnV5dGVI6P+iDpqykdt8iiwskN4GMNLj4Scrh8rjsC
R0SgqK96CwRsjeZoY7nEgLqCmN4hdDF7BxHqjcMzEzi896wesoJu40Yv4+Ei5LblAsyI2DAF+SyQ
iuk4gMuzimIYmZC5ROwui4XrKdlRpxoZBVM+aFhhluWeLmj3463yOvjZNrkCqn3I1CcaZZ8tUWDz
hxXpEGfbDXyo3dhnxn+3oMwW6tyXIKnIBSY546bYx/N54qG1QbQD9Vs1rABqlv5tkSKz6hNSl/ci
wuSNAV6z1Uiw5/RpV+dL+ah/RF0nkVRiga2VMfDVV7Abk79c8JGMqQShYil+kcK604MC/LQjwWZz
4FBDCVBZUgBujbJ6dXVbUkUOhecbKqQ1nW9cLEmR8ZvoVmTrcz8D7GccXgJFDRNy/h6GFSwtiXio
Ff2UhnnZYRTLBZFa5QMd5vVklvVI9pkS9LiIOJR77e22KhGujY6wZoHxtLgzpT7VxFo8hoMdp8Q+
Nv394tik+42eWoApv7cLhiastlGW/LSAhQJ1Gx4qiSDvIg5gMFm+TzVGTSSjAqBdtpkXs12vtP6K
OH1F/idMWkss4DUWiwOBmbMEBTFbthcvSX4uCbqsdoZVSmqF9HmZT9c6fHiRQ+5TOzvGRIdN7UCO
zqvqJzQ1c+SRq7Dnn6Cp9BlCxOGuk8rOa/PINUffb5bgs4BPpa1qX0K+XQDDRtcY5gZsSESu0sFP
+3eqtU+dZOYkGvBxPIQ/Lx3MqVllqwYs/MwXBV7JF9wlsAt471u4TN3Bj7iQ2S/KKbuGeIJk7AfF
oBIKMRKH9J6yU5kY72JooLDlSxfF2fTKGwmSLbwE6pjJ+EOxL0Ff4a/M24ocALp4/5AYXaBBqDKh
82qxYvsIv3CmZh6Ew0d92MTRrz1srsVsCFVwte6E9Y/Qf6PDcXplckxiEaM5pwwSENTFlL72evPR
CnRzxRCup/jyReWKah8ZVg7tyyO0YcOremT3P7ko2sJgaSNkinfaf5rNPKtl88AyGg9NBtZgW3Ph
szjsB33f/Mvdvlvfqw9KQ5oB7JXCBa6xg7ZsMDDnSnHzMNWaYOU4KsO5LRbmNDZxBp85HZnrq6Vq
WXI2fx0iRE1a6BuCXXq+BW3w1uNcHxB/2AiIYrJEY9oSmL+DWuW8k+aVirCSgYTYKFVO/n7PnUlN
o2Rnk2ibG0HWWn3Kau8ION9y2pk5+3Y8Bbcyf1kFUvtZfTC4k+Sa4M3JZ4namLAIplWSqQOsJQb2
SlZl9Ka5HTXBmqVcYxX/1wXKBXA13MRoQUDwjisKDChIEJzWgDPuiGIYr3aE5fR35FRS1TgNvLZx
4i1vAR2bWjbkTs69Zsml+RKoZ2vqiyig7djSO1lrRIyrmF8BMeU2Vy60NhMj+ZMpgfvF5hiJPLH7
c5M+vUbNTHd6WLXrRhXZhAQp9Zt27jIS0ltYZRc4as8MSoVopIQNIGAcNPiHigsZr0SvnmoY0qbP
P9IBj9D5Ax8zAFuVohetIY0OcxFvH3pM5L7MbL+0vPHERusZC1m1uJM8Xst+Xl2CiCbFY1mWeIBH
VPdH6K8YYggi/WYizrz0bT3mut+UZ1ClZSjNswx7EYZyTTJfmOpPAYHurHjm9nnSgyqPTh1nmus/
4YHTWxhcrcXJdRt3XEAxAHv3EVnAKYR16Zi6kDO2MyQp3U1oc0jWD3ofrVENo28wdv3B1CjrxiuY
Y4EZ2Ix5I/WH1KnjvGnUoPB1RAapObw2raV5YsIG4Sq1GIgDNcBRjzTIy27vlX/ANzfVwlxAVAcV
DWQ4X2umVUBbt+D3jxz0ODQkqXjEWYCgSFDCX4xiAjx7RCRFl7hXuqOMboA6x6vUWXZaZchnuSJw
kHFp/Ty/uOicermfvNzbJMMHeIOzUrMjS/wkqA2H6zhm59MZ3ERHXHdQExaGUrp0gMUyA6Fkcvse
dr0uQxYSE6LtGW6jetX6CAEA8+3rUCyS2mC5r0gWFwgzkoxZRFZVHfwCGfJ93+xrpnNDEJyIDc+K
o3SJIJYzsifIDIh6vxjJW+rYvj7D08q7r30bkmpYXouMzMajwg5TokmrJA78pPJg1AD1WEeRLl2s
msAx1WjMWMss0+prlbTMPLpJp1/5m/9+pSiPAo02Thac6mHnOGc3JeidEJLCrlrErff1pc7cdKbf
7/92Hmq/ZbO02UgvNjHAE7AH88F5B8mfkyrvdCuEUD2GTbzhfbKCn529s2t0NDXwKIcH5YPcwFyI
affJ71VhfkZsQ4pXy/THLtDAYOTGEIu6+LNgQ8mMOUdSl0UQR8GwqyAqkhR61Ub6LJNykV1m1ccv
6qyo//4v2BplZkKMo79EnytS+H0yigzwzGwm1v65oTlzIGDYzlJ5yCkfGzqcqI93uqSkFqRmwII8
l5ElK5iAt+ipd3Lt/2m519lDgkPnMjiHy94QsPFLMSjcNPlnlsOovFaBTWBDllzMN5RWLp9NayLg
l+irWY0WagtbqtZDsRrcnm37QCXKqmPg53qBgTY03OFpOCxoFMhY65mdyoCXXcoNgD7Hhav89kJz
NQszCA5LUIGmf1pjqa9R6l5NzaWAGN5HfzrWQOa7eIXlyE6H7nhbSqJbOB5M/GP7nTUOf67K6G2q
Qpb+1uYDbogThI7cbVEUruoA6zDYut5/q1LskR+60uGSnEmZK7OlD+m+Q+so6Yb+bQuLRsJ3whlM
NRpiLBIFZjLRhVxPfl3jIlkl2YKsEFi6S4REst5PkdipwSMbToaCpaUTYu00JNwq2x3tkH3GGv8u
XrB05cUgfHWDgaCPXJ9QbOEFjP9es1jDppuWmEZotKE4tUj3KXwBP37eK6quVMXzxyAyM+2THQdG
eY2gEVdjY2I39auwEE4K+TEun/Z8d1teJqxOD4JBfH5aGAvvDV832KsNmKFxdax/vvhtoKQ3O6W/
cjZjAi4Jn5Bz2zS11BcdZNEUrji4nqX+6vJ0K4siHK/R6bCS5+xKjKaDSsrlvhdK1D8Zh2lVBpip
1RlJ1fmIgvNOW4XskUwxBSCd1vrWExxoNjulc1WZ5jeCHDBccr4V0xEHic5Xaz8WHkZWkIfTRtF5
sRkG4WlMSDK71eUcZ1uMVUYQIwOwZerS/F3v/M5tluTzyC5wnF64XM72G62ZetoYwpki/d74fxGj
THiK9rQ4YMN8QqiPBBJLI2YPhi03wWVtegtLIg9yOfrEwK44SGzNswACHoXCkPWYOEbMUvmuAkMU
066MitNUTY3vfrLiWWjn/lKthUxsNh+nIx33BfyKAWcYGptuQ565OG30s6vD83vE28VTgXIR4UKR
iwvx+3U6C39vG9kBta+vFHbGrV0npcCiHjyU/6WuFfKivUMm6Lk0U9TPQHGjCa0+Q9vI8Qtg1ixD
GonUiKs4fcCU5QkXB06qrI2jx16mGS4CCy/yWMYbBbDIlPj++AvhI2KA7QmHugOEYQt6HyAzp+29
QdLrdBiZtmHDqUGoyMvT+wr8PI9ERxv1jAfR1xcVNr9Iq+Pw2nDg3H/LW7tPfVCRUcE6ZuZiVOJL
OXHQyc6gU6UD8LKDYxTM1sd42/V+juYu3FkFYoBrm3cP0San9e8b0nWjkMhj3ocXw5kYy6gpqXJi
VG0Ixf+jc5WCS90+AALU2t6BlUeScO87Sh4PHB5md94XmutjtjqTHikM26VhHy3YmGedl6AdngI=
`pragma protect end_protected
