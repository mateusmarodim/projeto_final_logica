-- system_0_lab7_final_0.vhd

-- Generated using ACDS version 13.0sp1 232 at 2024.07.03.21:10:14

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity system_0_lab7_final_0 is
	port (
		chipselect : in  std_logic                     := '0';             -- avalon_slave_0.chipselect
		writedata  : in  std_logic_vector(31 downto 0) := (others => '0'); --               .writedata
		readdata   : out std_logic_vector(31 downto 0);                    --               .readdata
		add        : in  std_logic                     := '0';             --               .address
		write_en   : in  std_logic                     := '0';             --               .write
		read_en    : in  std_logic                     := '0';             --               .read
		clock      : in  std_logic                     := '0';             --     clock_sink.clk
		resetn     : in  std_logic                     := '0'              --     reset_sink.reset_n
	);
end entity system_0_lab7_final_0;

architecture rtl of system_0_lab7_final_0 is
	component top_avalon is
		port (
			chipselect : in  std_logic                     := 'X';             -- chipselect
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			add        : in  std_logic                     := 'X';             -- address
			write_en   : in  std_logic                     := 'X';             -- write
			read_en    : in  std_logic                     := 'X';             -- read
			clock      : in  std_logic                     := 'X';             -- clk
			resetn     : in  std_logic                     := 'X'              -- reset_n
		);
	end component top_avalon;

begin

	lab7_final_0 : component top_avalon
		port map (
			chipselect => chipselect, -- avalon_slave_0.chipselect
			writedata  => writedata,  --               .writedata
			readdata   => readdata,   --               .readdata
			add        => add,        --               .address
			write_en   => write_en,   --               .write
			read_en    => read_en,    --               .read
			clock      => clock,      --     clock_sink.clk
			resetn     => resetn      --     reset_sink.reset_n
		);

end architecture rtl; -- of system_0_lab7_final_0
